
module weights_rom_depthwise_pointwise_2 (
    input wire [15:0] addr, 
    output reg [7:0] data) ;
    reg [7:0] rom [0:18431] ; 
    initial
        begin
            rom[0] = 8'hf3 ;
            rom[1] = 8'he7 ;
            rom[2] = 8'hf1 ;
            rom[3] = 8'h03 ;
            rom[4] = 8'h0a ;
            rom[5] = 8'h09 ;
            rom[6] = 8'hd8 ;
            rom[7] = 8'hb6 ;
            rom[8] = 8'hd8 ;
            rom[9] = 8'h11 ;
            rom[10] = 8'hfc ;
            rom[11] = 8'h0d ;
            rom[12] = 8'he5 ;
            rom[13] = 8'hd8 ;
            rom[14] = 8'h23 ;
            rom[15] = 8'h15 ;
            rom[16] = 8'hec ;
            rom[17] = 8'hef ;
            rom[18] = 8'h06 ;
            rom[19] = 8'hf6 ;
            rom[20] = 8'hf8 ;
            rom[21] = 8'h05 ;
            rom[22] = 8'h0d ;
            rom[23] = 8'hf0 ;
            rom[24] = 8'hda ;
            rom[25] = 8'h07 ;
            rom[26] = 8'hf6 ;
            rom[27] = 8'h05 ;
            rom[28] = 8'hfc ;
            rom[29] = 8'hde ;
            rom[30] = 8'hee ;
            rom[31] = 8'h03 ;
            rom[32] = 8'hfd ;
            rom[33] = 8'he1 ;
            rom[34] = 8'h08 ;
            rom[35] = 8'hfa ;
            rom[36] = 8'hdb ;
            rom[37] = 8'hf4 ;
            rom[38] = 8'h1a ;
            rom[39] = 8'hfb ;
            rom[40] = 8'hf3 ;
            rom[41] = 8'hee ;
            rom[42] = 8'hcd ;
            rom[43] = 8'hfb ;
            rom[44] = 8'h09 ;
            rom[45] = 8'hf9 ;
            rom[46] = 8'h19 ;
            rom[47] = 8'hf2 ;
            rom[48] = 8'hec ;
            rom[49] = 8'h17 ;
            rom[50] = 8'hef ;
            rom[51] = 8'h18 ;
            rom[52] = 8'hf0 ;
            rom[53] = 8'hea ;
            rom[54] = 8'h06 ;
            rom[55] = 8'he7 ;
            rom[56] = 8'h11 ;
            rom[57] = 8'h14 ;
            rom[58] = 8'hc0 ;
            rom[59] = 8'hd6 ;
            rom[60] = 8'h04 ;
            rom[61] = 8'h09 ;
            rom[62] = 8'h11 ;
            rom[63] = 8'hf7 ;
            rom[64] = 8'h17 ;
            rom[65] = 8'h09 ;
            rom[66] = 8'h0d ;
            rom[67] = 8'h01 ;
            rom[68] = 8'h17 ;
            rom[69] = 8'hfe ;
            rom[70] = 8'he4 ;
            rom[71] = 8'h09 ;
            rom[72] = 8'hf6 ;
            rom[73] = 8'h06 ;
            rom[74] = 8'hf2 ;
            rom[75] = 8'h06 ;
            rom[76] = 8'h0c ;
            rom[77] = 8'hf7 ;
            rom[78] = 8'hfa ;
            rom[79] = 8'h10 ;
            rom[80] = 8'hf9 ;
            rom[81] = 8'h0b ;
            rom[82] = 8'hd8 ;
            rom[83] = 8'h1a ;
            rom[84] = 8'hf6 ;
            rom[85] = 8'h18 ;
            rom[86] = 8'hfe ;
            rom[87] = 8'h01 ;
            rom[88] = 8'h10 ;
            rom[89] = 8'h11 ;
            rom[90] = 8'h02 ;
            rom[91] = 8'hf7 ;
            rom[92] = 8'h0d ;
            rom[93] = 8'hf0 ;
            rom[94] = 8'h1d ;
            rom[95] = 8'he4 ;
            rom[96] = 8'h0f ;
            rom[97] = 8'hee ;
            rom[98] = 8'hd1 ;
            rom[99] = 8'h13 ;
            rom[100] = 8'h12 ;
            rom[101] = 8'hf7 ;
            rom[102] = 8'hf9 ;
            rom[103] = 8'h00 ;
            rom[104] = 8'h06 ;
            rom[105] = 8'hfc ;
            rom[106] = 8'hf5 ;
            rom[107] = 8'h20 ;
            rom[108] = 8'h05 ;
            rom[109] = 8'h0e ;
            rom[110] = 8'h20 ;
            rom[111] = 8'h09 ;
            rom[112] = 8'h12 ;
            rom[113] = 8'h03 ;
            rom[114] = 8'h06 ;
            rom[115] = 8'h09 ;
            rom[116] = 8'h07 ;
            rom[117] = 8'h0a ;
            rom[118] = 8'h11 ;
            rom[119] = 8'hea ;
            rom[120] = 8'h20 ;
            rom[121] = 8'hff ;
            rom[122] = 8'hd0 ;
            rom[123] = 8'h06 ;
            rom[124] = 8'h0f ;
            rom[125] = 8'hec ;
            rom[126] = 8'h24 ;
            rom[127] = 8'h05 ;
            rom[128] = 8'hff ;
            rom[129] = 8'he5 ;
            rom[130] = 8'h06 ;
            rom[131] = 8'h18 ;
            rom[132] = 8'h13 ;
            rom[133] = 8'hfa ;
            rom[134] = 8'hef ;
            rom[135] = 8'h1e ;
            rom[136] = 8'h00 ;
            rom[137] = 8'hf3 ;
            rom[138] = 8'hf8 ;
            rom[139] = 8'h01 ;
            rom[140] = 8'hf2 ;
            rom[141] = 8'hed ;
            rom[142] = 8'h16 ;
            rom[143] = 8'hfd ;
            rom[144] = 8'hf6 ;
            rom[145] = 8'h07 ;
            rom[146] = 8'hd8 ;
            rom[147] = 8'h0e ;
            rom[148] = 8'h03 ;
            rom[149] = 8'he4 ;
            rom[150] = 8'h0d ;
            rom[151] = 8'hff ;
            rom[152] = 8'hfc ;
            rom[153] = 8'h08 ;
            rom[154] = 8'h0c ;
            rom[155] = 8'h0e ;
            rom[156] = 8'hf3 ;
            rom[157] = 8'hf0 ;
            rom[158] = 8'h1b ;
            rom[159] = 8'hf3 ;
            rom[160] = 8'hfa ;
            rom[161] = 8'he2 ;
            rom[162] = 8'h17 ;
            rom[163] = 8'hf3 ;
            rom[164] = 8'hf3 ;
            rom[165] = 8'hf6 ;
            rom[166] = 8'he4 ;
            rom[167] = 8'hfc ;
            rom[168] = 8'hea ;
            rom[169] = 8'hf3 ;
            rom[170] = 8'hf5 ;
            rom[171] = 8'h04 ;
            rom[172] = 8'hf2 ;
            rom[173] = 8'h28 ;
            rom[174] = 8'hed ;
            rom[175] = 8'h0f ;
            rom[176] = 8'hfc ;
            rom[177] = 8'h1d ;
            rom[178] = 8'h11 ;
            rom[179] = 8'h14 ;
            rom[180] = 8'hff ;
            rom[181] = 8'hd3 ;
            rom[182] = 8'hfa ;
            rom[183] = 8'h0d ;
            rom[184] = 8'he5 ;
            rom[185] = 8'hec ;
            rom[186] = 8'h01 ;
            rom[187] = 8'h07 ;
            rom[188] = 8'hd0 ;
            rom[189] = 8'hfd ;
            rom[190] = 8'h1d ;
            rom[191] = 8'hf9 ;
            rom[192] = 8'hf4 ;
            rom[193] = 8'h06 ;
            rom[194] = 8'hdd ;
            rom[195] = 8'h35 ;
            rom[196] = 8'h18 ;
            rom[197] = 8'h1b ;
            rom[198] = 8'hc2 ;
            rom[199] = 8'hf7 ;
            rom[200] = 8'h1f ;
            rom[201] = 8'hec ;
            rom[202] = 8'hed ;
            rom[203] = 8'h01 ;
            rom[204] = 8'h08 ;
            rom[205] = 8'hf7 ;
            rom[206] = 8'h19 ;
            rom[207] = 8'hf8 ;
            rom[208] = 8'hff ;
            rom[209] = 8'h12 ;
            rom[210] = 8'hff ;
            rom[211] = 8'he9 ;
            rom[212] = 8'hf7 ;
            rom[213] = 8'h06 ;
            rom[214] = 8'h08 ;
            rom[215] = 8'hdc ;
            rom[216] = 8'h02 ;
            rom[217] = 8'h20 ;
            rom[218] = 8'hf3 ;
            rom[219] = 8'he9 ;
            rom[220] = 8'he6 ;
            rom[221] = 8'hee ;
            rom[222] = 8'h10 ;
            rom[223] = 8'h11 ;
            rom[224] = 8'hff ;
            rom[225] = 8'h11 ;
            rom[226] = 8'h18 ;
            rom[227] = 8'h1d ;
            rom[228] = 8'h17 ;
            rom[229] = 8'hfe ;
            rom[230] = 8'h05 ;
            rom[231] = 8'he5 ;
            rom[232] = 8'he7 ;
            rom[233] = 8'hfb ;
            rom[234] = 8'hdb ;
            rom[235] = 8'h22 ;
            rom[236] = 8'h20 ;
            rom[237] = 8'hf8 ;
            rom[238] = 8'h01 ;
            rom[239] = 8'hf2 ;
            rom[240] = 8'h06 ;
            rom[241] = 8'hf8 ;
            rom[242] = 8'h0c ;
            rom[243] = 8'h02 ;
            rom[244] = 8'hdd ;
            rom[245] = 8'hed ;
            rom[246] = 8'he9 ;
            rom[247] = 8'h0b ;
            rom[248] = 8'hf6 ;
            rom[249] = 8'hfc ;
            rom[250] = 8'h12 ;
            rom[251] = 8'h13 ;
            rom[252] = 8'hcd ;
            rom[253] = 8'h0a ;
            rom[254] = 8'h04 ;
            rom[255] = 8'h0c ;
            rom[256] = 8'h19 ;
            rom[257] = 8'hf8 ;
            rom[258] = 8'hf5 ;
            rom[259] = 8'hef ;
            rom[260] = 8'h19 ;
            rom[261] = 8'h03 ;
            rom[262] = 8'h06 ;
            rom[263] = 8'h0e ;
            rom[264] = 8'hfb ;
            rom[265] = 8'h02 ;
            rom[266] = 8'he7 ;
            rom[267] = 8'he1 ;
            rom[268] = 8'h0d ;
            rom[269] = 8'h04 ;
            rom[270] = 8'hf6 ;
            rom[271] = 8'h1a ;
            rom[272] = 8'h08 ;
            rom[273] = 8'hf9 ;
            rom[274] = 8'hed ;
            rom[275] = 8'h03 ;
            rom[276] = 8'h0d ;
            rom[277] = 8'hd4 ;
            rom[278] = 8'h0b ;
            rom[279] = 8'h10 ;
            rom[280] = 8'h1c ;
            rom[281] = 8'h0d ;
            rom[282] = 8'he4 ;
            rom[283] = 8'h18 ;
            rom[284] = 8'h13 ;
            rom[285] = 8'hfa ;
            rom[286] = 8'h0a ;
            rom[287] = 8'hed ;
            rom[288] = 8'h06 ;
            rom[289] = 8'h09 ;
            rom[290] = 8'hfc ;
            rom[291] = 8'hcf ;
            rom[292] = 8'h09 ;
            rom[293] = 8'h14 ;
            rom[294] = 8'h07 ;
            rom[295] = 8'hf8 ;
            rom[296] = 8'hf2 ;
            rom[297] = 8'hbd ;
            rom[298] = 8'hff ;
            rom[299] = 8'hfa ;
            rom[300] = 8'h01 ;
            rom[301] = 8'h13 ;
            rom[302] = 8'hec ;
            rom[303] = 8'h01 ;
            rom[304] = 8'he4 ;
            rom[305] = 8'h2d ;
            rom[306] = 8'hf0 ;
            rom[307] = 8'he2 ;
            rom[308] = 8'hfc ;
            rom[309] = 8'he4 ;
            rom[310] = 8'hf6 ;
            rom[311] = 8'hf6 ;
            rom[312] = 8'hfa ;
            rom[313] = 8'hf6 ;
            rom[314] = 8'hfb ;
            rom[315] = 8'h0c ;
            rom[316] = 8'h0d ;
            rom[317] = 8'h10 ;
            rom[318] = 8'he0 ;
            rom[319] = 8'h09 ;
            rom[320] = 8'h09 ;
            rom[321] = 8'h1d ;
            rom[322] = 8'he6 ;
            rom[323] = 8'hfa ;
            rom[324] = 8'hfc ;
            rom[325] = 8'hf2 ;
            rom[326] = 8'hfd ;
            rom[327] = 8'h05 ;
            rom[328] = 8'h05 ;
            rom[329] = 8'he0 ;
            rom[330] = 8'h05 ;
            rom[331] = 8'h14 ;
            rom[332] = 8'h0c ;
            rom[333] = 8'hed ;
            rom[334] = 8'hee ;
            rom[335] = 8'h11 ;
            rom[336] = 8'h10 ;
            rom[337] = 8'h09 ;
            rom[338] = 8'hf1 ;
            rom[339] = 8'hfd ;
            rom[340] = 8'hfc ;
            rom[341] = 8'h17 ;
            rom[342] = 8'heb ;
            rom[343] = 8'h03 ;
            rom[344] = 8'hf9 ;
            rom[345] = 8'h29 ;
            rom[346] = 8'he3 ;
            rom[347] = 8'h06 ;
            rom[348] = 8'hf4 ;
            rom[349] = 8'h20 ;
            rom[350] = 8'hfb ;
            rom[351] = 8'h18 ;
            rom[352] = 8'hef ;
            rom[353] = 8'h17 ;
            rom[354] = 8'hd3 ;
            rom[355] = 8'hfa ;
            rom[356] = 8'h15 ;
            rom[357] = 8'hea ;
            rom[358] = 8'hd3 ;
            rom[359] = 8'h12 ;
            rom[360] = 8'hf5 ;
            rom[361] = 8'h03 ;
            rom[362] = 8'h01 ;
            rom[363] = 8'hce ;
            rom[364] = 8'hea ;
            rom[365] = 8'h01 ;
            rom[366] = 8'h19 ;
            rom[367] = 8'hfb ;
            rom[368] = 8'h07 ;
            rom[369] = 8'hf4 ;
            rom[370] = 8'h09 ;
            rom[371] = 8'heb ;
            rom[372] = 8'he0 ;
            rom[373] = 8'h0f ;
            rom[374] = 8'h10 ;
            rom[375] = 8'h1a ;
            rom[376] = 8'hf0 ;
            rom[377] = 8'hf3 ;
            rom[378] = 8'h16 ;
            rom[379] = 8'h05 ;
            rom[380] = 8'hf7 ;
            rom[381] = 8'hf4 ;
            rom[382] = 8'hf8 ;
            rom[383] = 8'hf8 ;
            rom[384] = 8'h08 ;
            rom[385] = 8'hf0 ;
            rom[386] = 8'hef ;
            rom[387] = 8'hfc ;
            rom[388] = 8'h06 ;
            rom[389] = 8'h0d ;
            rom[390] = 8'h0c ;
            rom[391] = 8'hfc ;
            rom[392] = 8'he7 ;
            rom[393] = 8'hf5 ;
            rom[394] = 8'h0a ;
            rom[395] = 8'hfd ;
            rom[396] = 8'h09 ;
            rom[397] = 8'hf0 ;
            rom[398] = 8'h08 ;
            rom[399] = 8'h07 ;
            rom[400] = 8'h01 ;
            rom[401] = 8'hf0 ;
            rom[402] = 8'h0c ;
            rom[403] = 8'hf9 ;
            rom[404] = 8'h00 ;
            rom[405] = 8'h12 ;
            rom[406] = 8'h1e ;
            rom[407] = 8'he8 ;
            rom[408] = 8'hd5 ;
            rom[409] = 8'h13 ;
            rom[410] = 8'h0f ;
            rom[411] = 8'h0a ;
            rom[412] = 8'hff ;
            rom[413] = 8'hf3 ;
            rom[414] = 8'h17 ;
            rom[415] = 8'he9 ;
            rom[416] = 8'hef ;
            rom[417] = 8'hf0 ;
            rom[418] = 8'h17 ;
            rom[419] = 8'hd0 ;
            rom[420] = 8'hf8 ;
            rom[421] = 8'h0a ;
            rom[422] = 8'h0d ;
            rom[423] = 8'hf7 ;
            rom[424] = 8'hf5 ;
            rom[425] = 8'h13 ;
            rom[426] = 8'he9 ;
            rom[427] = 8'hf4 ;
            rom[428] = 8'h20 ;
            rom[429] = 8'hf8 ;
            rom[430] = 8'h0d ;
            rom[431] = 8'hfb ;
            rom[432] = 8'h0d ;
            rom[433] = 8'h17 ;
            rom[434] = 8'hd2 ;
            rom[435] = 8'hff ;
            rom[436] = 8'h09 ;
            rom[437] = 8'h07 ;
            rom[438] = 8'h0c ;
            rom[439] = 8'h2c ;
            rom[440] = 8'hec ;
            rom[441] = 8'h1b ;
            rom[442] = 8'hdf ;
            rom[443] = 8'h2e ;
            rom[444] = 8'hd2 ;
            rom[445] = 8'hd7 ;
            rom[446] = 8'h14 ;
            rom[447] = 8'h08 ;
            rom[448] = 8'heb ;
            rom[449] = 8'hc4 ;
            rom[450] = 8'h02 ;
            rom[451] = 8'hfd ;
            rom[452] = 8'h08 ;
            rom[453] = 8'h08 ;
            rom[454] = 8'hd6 ;
            rom[455] = 8'hf1 ;
            rom[456] = 8'he9 ;
            rom[457] = 8'hf3 ;
            rom[458] = 8'h0a ;
            rom[459] = 8'h04 ;
            rom[460] = 8'h1f ;
            rom[461] = 8'he9 ;
            rom[462] = 8'h08 ;
            rom[463] = 8'he2 ;
            rom[464] = 8'h04 ;
            rom[465] = 8'h00 ;
            rom[466] = 8'he0 ;
            rom[467] = 8'he6 ;
            rom[468] = 8'h09 ;
            rom[469] = 8'he3 ;
            rom[470] = 8'hf0 ;
            rom[471] = 8'h0d ;
            rom[472] = 8'h16 ;
            rom[473] = 8'h02 ;
            rom[474] = 8'h08 ;
            rom[475] = 8'he3 ;
            rom[476] = 8'h2e ;
            rom[477] = 8'hdc ;
            rom[478] = 8'h00 ;
            rom[479] = 8'h23 ;
            rom[480] = 8'h11 ;
            rom[481] = 8'h04 ;
            rom[482] = 8'h04 ;
            rom[483] = 8'h2a ;
            rom[484] = 8'h25 ;
            rom[485] = 8'h16 ;
            rom[486] = 8'hed ;
            rom[487] = 8'h02 ;
            rom[488] = 8'hfc ;
            rom[489] = 8'h03 ;
            rom[490] = 8'hd9 ;
            rom[491] = 8'h11 ;
            rom[492] = 8'h0f ;
            rom[493] = 8'h09 ;
            rom[494] = 8'h09 ;
            rom[495] = 8'h28 ;
            rom[496] = 8'h0d ;
            rom[497] = 8'hfc ;
            rom[498] = 8'h12 ;
            rom[499] = 8'h06 ;
            rom[500] = 8'hdd ;
            rom[501] = 8'he5 ;
            rom[502] = 8'h0d ;
            rom[503] = 8'h00 ;
            rom[504] = 8'h00 ;
            rom[505] = 8'hf9 ;
            rom[506] = 8'hf1 ;
            rom[507] = 8'h0d ;
            rom[508] = 8'hda ;
            rom[509] = 8'hdd ;
            rom[510] = 8'h30 ;
            rom[511] = 8'h00 ;
            rom[512] = 8'hec ;
            rom[513] = 8'h2b ;
            rom[514] = 8'h16 ;
            rom[515] = 8'hec ;
            rom[516] = 8'h0b ;
            rom[517] = 8'h11 ;
            rom[518] = 8'h01 ;
            rom[519] = 8'h14 ;
            rom[520] = 8'hff ;
            rom[521] = 8'hf8 ;
            rom[522] = 8'hf4 ;
            rom[523] = 8'h04 ;
            rom[524] = 8'he5 ;
            rom[525] = 8'hfd ;
            rom[526] = 8'h0c ;
            rom[527] = 8'h11 ;
            rom[528] = 8'h0e ;
            rom[529] = 8'h0f ;
            rom[530] = 8'hff ;
            rom[531] = 8'hfd ;
            rom[532] = 8'h01 ;
            rom[533] = 8'h0f ;
            rom[534] = 8'hf9 ;
            rom[535] = 8'hf8 ;
            rom[536] = 8'h15 ;
            rom[537] = 8'h04 ;
            rom[538] = 8'h02 ;
            rom[539] = 8'hed ;
            rom[540] = 8'h15 ;
            rom[541] = 8'hfe ;
            rom[542] = 8'hfe ;
            rom[543] = 8'hca ;
            rom[544] = 8'hff ;
            rom[545] = 8'hf9 ;
            rom[546] = 8'hdd ;
            rom[547] = 8'h1c ;
            rom[548] = 8'h0e ;
            rom[549] = 8'hea ;
            rom[550] = 8'heb ;
            rom[551] = 8'heb ;
            rom[552] = 8'h0e ;
            rom[553] = 8'hd0 ;
            rom[554] = 8'h16 ;
            rom[555] = 8'hf4 ;
            rom[556] = 8'h00 ;
            rom[557] = 8'hff ;
            rom[558] = 8'hf1 ;
            rom[559] = 8'h09 ;
            rom[560] = 8'h01 ;
            rom[561] = 8'hdf ;
            rom[562] = 8'h02 ;
            rom[563] = 8'he0 ;
            rom[564] = 8'h12 ;
            rom[565] = 8'h0f ;
            rom[566] = 8'hf4 ;
            rom[567] = 8'h0f ;
            rom[568] = 8'hf0 ;
            rom[569] = 8'hfe ;
            rom[570] = 8'hf6 ;
            rom[571] = 8'h14 ;
            rom[572] = 8'h06 ;
            rom[573] = 8'h17 ;
            rom[574] = 8'h08 ;
            rom[575] = 8'h13 ;
            rom[576] = 8'h1c ;
            rom[577] = 8'h11 ;
            rom[578] = 8'h1f ;
            rom[579] = 8'hd8 ;
            rom[580] = 8'h04 ;
            rom[581] = 8'h02 ;
            rom[582] = 8'h04 ;
            rom[583] = 8'h05 ;
            rom[584] = 8'hfe ;
            rom[585] = 8'h1b ;
            rom[586] = 8'h0d ;
            rom[587] = 8'he8 ;
            rom[588] = 8'hf2 ;
            rom[589] = 8'he9 ;
            rom[590] = 8'h03 ;
            rom[591] = 8'h04 ;
            rom[592] = 8'hfb ;
            rom[593] = 8'h05 ;
            rom[594] = 8'hfc ;
            rom[595] = 8'h05 ;
            rom[596] = 8'hee ;
            rom[597] = 8'heb ;
            rom[598] = 8'hfc ;
            rom[599] = 8'h0f ;
            rom[600] = 8'hfd ;
            rom[601] = 8'hf1 ;
            rom[602] = 8'hf7 ;
            rom[603] = 8'hed ;
            rom[604] = 8'h09 ;
            rom[605] = 8'h06 ;
            rom[606] = 8'hf8 ;
            rom[607] = 8'hbc ;
            rom[608] = 8'hef ;
            rom[609] = 8'h01 ;
            rom[610] = 8'he7 ;
            rom[611] = 8'h10 ;
            rom[612] = 8'h13 ;
            rom[613] = 8'he5 ;
            rom[614] = 8'h02 ;
            rom[615] = 8'he7 ;
            rom[616] = 8'h0c ;
            rom[617] = 8'he5 ;
            rom[618] = 8'h0b ;
            rom[619] = 8'h05 ;
            rom[620] = 8'hdf ;
            rom[621] = 8'h01 ;
            rom[622] = 8'hfd ;
            rom[623] = 8'h0c ;
            rom[624] = 8'h1a ;
            rom[625] = 8'hf2 ;
            rom[626] = 8'he0 ;
            rom[627] = 8'hfc ;
            rom[628] = 8'h0d ;
            rom[629] = 8'hef ;
            rom[630] = 8'h05 ;
            rom[631] = 8'h12 ;
            rom[632] = 8'hdc ;
            rom[633] = 8'h05 ;
            rom[634] = 8'heb ;
            rom[635] = 8'h12 ;
            rom[636] = 8'hff ;
            rom[637] = 8'hf3 ;
            rom[638] = 8'h00 ;
            rom[639] = 8'h01 ;
            rom[640] = 8'he5 ;
            rom[641] = 8'h07 ;
            rom[642] = 8'he7 ;
            rom[643] = 8'hf8 ;
            rom[644] = 8'h13 ;
            rom[645] = 8'h08 ;
            rom[646] = 8'hfe ;
            rom[647] = 8'he4 ;
            rom[648] = 8'h05 ;
            rom[649] = 8'hf7 ;
            rom[650] = 8'h16 ;
            rom[651] = 8'h07 ;
            rom[652] = 8'h09 ;
            rom[653] = 8'h02 ;
            rom[654] = 8'h0a ;
            rom[655] = 8'hfb ;
            rom[656] = 8'h17 ;
            rom[657] = 8'h04 ;
            rom[658] = 8'hda ;
            rom[659] = 8'h1c ;
            rom[660] = 8'h05 ;
            rom[661] = 8'h26 ;
            rom[662] = 8'hd5 ;
            rom[663] = 8'hfa ;
            rom[664] = 8'h19 ;
            rom[665] = 8'hf7 ;
            rom[666] = 8'hf2 ;
            rom[667] = 8'hc7 ;
            rom[668] = 8'h0c ;
            rom[669] = 8'h19 ;
            rom[670] = 8'h2b ;
            rom[671] = 8'hf0 ;
            rom[672] = 8'h06 ;
            rom[673] = 8'h11 ;
            rom[674] = 8'h1a ;
            rom[675] = 8'hf6 ;
            rom[676] = 8'hf1 ;
            rom[677] = 8'hf3 ;
            rom[678] = 8'hef ;
            rom[679] = 8'hfa ;
            rom[680] = 8'h0a ;
            rom[681] = 8'hfb ;
            rom[682] = 8'h00 ;
            rom[683] = 8'hf8 ;
            rom[684] = 8'h0f ;
            rom[685] = 8'hfd ;
            rom[686] = 8'h0b ;
            rom[687] = 8'hf9 ;
            rom[688] = 8'hea ;
            rom[689] = 8'h15 ;
            rom[690] = 8'h0b ;
            rom[691] = 8'h1c ;
            rom[692] = 8'hd6 ;
            rom[693] = 8'hff ;
            rom[694] = 8'h14 ;
            rom[695] = 8'he8 ;
            rom[696] = 8'h14 ;
            rom[697] = 8'h1b ;
            rom[698] = 8'he7 ;
            rom[699] = 8'h1f ;
            rom[700] = 8'h08 ;
            rom[701] = 8'he9 ;
            rom[702] = 8'hfc ;
            rom[703] = 8'hf4 ;
            rom[704] = 8'h18 ;
            rom[705] = 8'h29 ;
            rom[706] = 8'hff ;
            rom[707] = 8'h15 ;
            rom[708] = 8'h03 ;
            rom[709] = 8'h13 ;
            rom[710] = 8'h01 ;
            rom[711] = 8'hea ;
            rom[712] = 8'h05 ;
            rom[713] = 8'hde ;
            rom[714] = 8'hfa ;
            rom[715] = 8'h0f ;
            rom[716] = 8'h19 ;
            rom[717] = 8'h02 ;
            rom[718] = 8'h15 ;
            rom[719] = 8'hfd ;
            rom[720] = 8'h13 ;
            rom[721] = 8'h27 ;
            rom[722] = 8'h09 ;
            rom[723] = 8'hdd ;
            rom[724] = 8'hf7 ;
            rom[725] = 8'h0e ;
            rom[726] = 8'hfe ;
            rom[727] = 8'hf5 ;
            rom[728] = 8'he4 ;
            rom[729] = 8'h0a ;
            rom[730] = 8'h09 ;
            rom[731] = 8'h06 ;
            rom[732] = 8'h03 ;
            rom[733] = 8'h06 ;
            rom[734] = 8'h0a ;
            rom[735] = 8'h01 ;
            rom[736] = 8'h04 ;
            rom[737] = 8'h0f ;
            rom[738] = 8'h02 ;
            rom[739] = 8'h11 ;
            rom[740] = 8'hde ;
            rom[741] = 8'h09 ;
            rom[742] = 8'hee ;
            rom[743] = 8'hf3 ;
            rom[744] = 8'hf1 ;
            rom[745] = 8'hff ;
            rom[746] = 8'h20 ;
            rom[747] = 8'he1 ;
            rom[748] = 8'h22 ;
            rom[749] = 8'h21 ;
            rom[750] = 8'he5 ;
            rom[751] = 8'hf8 ;
            rom[752] = 8'h1e ;
            rom[753] = 8'h12 ;
            rom[754] = 8'h01 ;
            rom[755] = 8'h07 ;
            rom[756] = 8'h0d ;
            rom[757] = 8'h0a ;
            rom[758] = 8'h14 ;
            rom[759] = 8'hdb ;
            rom[760] = 8'h00 ;
            rom[761] = 8'h04 ;
            rom[762] = 8'hfc ;
            rom[763] = 8'hf5 ;
            rom[764] = 8'hf4 ;
            rom[765] = 8'h29 ;
            rom[766] = 8'h14 ;
            rom[767] = 8'h08 ;
            rom[768] = 8'hf8 ;
            rom[769] = 8'hf5 ;
            rom[770] = 8'h0c ;
            rom[771] = 8'h12 ;
            rom[772] = 8'hfc ;
            rom[773] = 8'h06 ;
            rom[774] = 8'he7 ;
            rom[775] = 8'h19 ;
            rom[776] = 8'hd0 ;
            rom[777] = 8'h0e ;
            rom[778] = 8'hee ;
            rom[779] = 8'h1a ;
            rom[780] = 8'h07 ;
            rom[781] = 8'hfc ;
            rom[782] = 8'h10 ;
            rom[783] = 8'h1c ;
            rom[784] = 8'hf5 ;
            rom[785] = 8'he2 ;
            rom[786] = 8'h09 ;
            rom[787] = 8'h00 ;
            rom[788] = 8'hf3 ;
            rom[789] = 8'h03 ;
            rom[790] = 8'hf5 ;
            rom[791] = 8'h17 ;
            rom[792] = 8'hf2 ;
            rom[793] = 8'h09 ;
            rom[794] = 8'h17 ;
            rom[795] = 8'he7 ;
            rom[796] = 8'hed ;
            rom[797] = 8'hfa ;
            rom[798] = 8'h17 ;
            rom[799] = 8'h10 ;
            rom[800] = 8'hf2 ;
            rom[801] = 8'hd9 ;
            rom[802] = 8'hfd ;
            rom[803] = 8'he7 ;
            rom[804] = 8'h04 ;
            rom[805] = 8'hfb ;
            rom[806] = 8'h0e ;
            rom[807] = 8'hed ;
            rom[808] = 8'h0b ;
            rom[809] = 8'hf5 ;
            rom[810] = 8'hda ;
            rom[811] = 8'h1d ;
            rom[812] = 8'h16 ;
            rom[813] = 8'h2a ;
            rom[814] = 8'h04 ;
            rom[815] = 8'h15 ;
            rom[816] = 8'hf4 ;
            rom[817] = 8'hfa ;
            rom[818] = 8'he0 ;
            rom[819] = 8'h13 ;
            rom[820] = 8'h04 ;
            rom[821] = 8'hed ;
            rom[822] = 8'h0c ;
            rom[823] = 8'h00 ;
            rom[824] = 8'h05 ;
            rom[825] = 8'h1a ;
            rom[826] = 8'hcc ;
            rom[827] = 8'h2a ;
            rom[828] = 8'he2 ;
            rom[829] = 8'hdc ;
            rom[830] = 8'h07 ;
            rom[831] = 8'h16 ;
            rom[832] = 8'h01 ;
            rom[833] = 8'h08 ;
            rom[834] = 8'h04 ;
            rom[835] = 8'h09 ;
            rom[836] = 8'hfb ;
            rom[837] = 8'h09 ;
            rom[838] = 8'hd7 ;
            rom[839] = 8'hf0 ;
            rom[840] = 8'hdb ;
            rom[841] = 8'hfe ;
            rom[842] = 8'h0d ;
            rom[843] = 8'hf6 ;
            rom[844] = 8'he1 ;
            rom[845] = 8'heb ;
            rom[846] = 8'hfe ;
            rom[847] = 8'h18 ;
            rom[848] = 8'h10 ;
            rom[849] = 8'hfa ;
            rom[850] = 8'h0d ;
            rom[851] = 8'hbf ;
            rom[852] = 8'hf9 ;
            rom[853] = 8'hf4 ;
            rom[854] = 8'h05 ;
            rom[855] = 8'h1a ;
            rom[856] = 8'hfd ;
            rom[857] = 8'h15 ;
            rom[858] = 8'he2 ;
            rom[859] = 8'hfb ;
            rom[860] = 8'h00 ;
            rom[861] = 8'h13 ;
            rom[862] = 8'h0c ;
            rom[863] = 8'h26 ;
            rom[864] = 8'hed ;
            rom[865] = 8'h0f ;
            rom[866] = 8'hf0 ;
            rom[867] = 8'h03 ;
            rom[868] = 8'h0b ;
            rom[869] = 8'hf6 ;
            rom[870] = 8'h25 ;
            rom[871] = 8'h08 ;
            rom[872] = 8'hf3 ;
            rom[873] = 8'h13 ;
            rom[874] = 8'hfb ;
            rom[875] = 8'hf2 ;
            rom[876] = 8'hfd ;
            rom[877] = 8'h3a ;
            rom[878] = 8'hf5 ;
            rom[879] = 8'h07 ;
            rom[880] = 8'hf9 ;
            rom[881] = 8'h03 ;
            rom[882] = 8'hf4 ;
            rom[883] = 8'hf0 ;
            rom[884] = 8'h01 ;
            rom[885] = 8'h02 ;
            rom[886] = 8'hfc ;
            rom[887] = 8'h1b ;
            rom[888] = 8'h00 ;
            rom[889] = 8'h0d ;
            rom[890] = 8'hdc ;
            rom[891] = 8'hfb ;
            rom[892] = 8'hdb ;
            rom[893] = 8'h22 ;
            rom[894] = 8'hf1 ;
            rom[895] = 8'h2c ;
            rom[896] = 8'h04 ;
            rom[897] = 8'h02 ;
            rom[898] = 8'h1b ;
            rom[899] = 8'h1e ;
            rom[900] = 8'h11 ;
            rom[901] = 8'h04 ;
            rom[902] = 8'he4 ;
            rom[903] = 8'h04 ;
            rom[904] = 8'hf0 ;
            rom[905] = 8'h01 ;
            rom[906] = 8'h02 ;
            rom[907] = 8'h11 ;
            rom[908] = 8'h03 ;
            rom[909] = 8'he6 ;
            rom[910] = 8'h04 ;
            rom[911] = 8'h0b ;
            rom[912] = 8'h00 ;
            rom[913] = 8'hf3 ;
            rom[914] = 8'h1a ;
            rom[915] = 8'hdc ;
            rom[916] = 8'he3 ;
            rom[917] = 8'h25 ;
            rom[918] = 8'h24 ;
            rom[919] = 8'hff ;
            rom[920] = 8'hed ;
            rom[921] = 8'hee ;
            rom[922] = 8'heb ;
            rom[923] = 8'hf8 ;
            rom[924] = 8'hfe ;
            rom[925] = 8'h06 ;
            rom[926] = 8'h12 ;
            rom[927] = 8'he1 ;
            rom[928] = 8'h0f ;
            rom[929] = 8'hf0 ;
            rom[930] = 8'h19 ;
            rom[931] = 8'h1a ;
            rom[932] = 8'hf7 ;
            rom[933] = 8'he6 ;
            rom[934] = 8'h02 ;
            rom[935] = 8'h08 ;
            rom[936] = 8'hda ;
            rom[937] = 8'h09 ;
            rom[938] = 8'hec ;
            rom[939] = 8'hff ;
            rom[940] = 8'hd5 ;
            rom[941] = 8'h17 ;
            rom[942] = 8'h17 ;
            rom[943] = 8'hd5 ;
            rom[944] = 8'h22 ;
            rom[945] = 8'h09 ;
            rom[946] = 8'hf0 ;
            rom[947] = 8'h11 ;
            rom[948] = 8'hee ;
            rom[949] = 8'h03 ;
            rom[950] = 8'h0f ;
            rom[951] = 8'hfc ;
            rom[952] = 8'h04 ;
            rom[953] = 8'hfa ;
            rom[954] = 8'hf9 ;
            rom[955] = 8'hf5 ;
            rom[956] = 8'h03 ;
            rom[957] = 8'hf5 ;
            rom[958] = 8'h02 ;
            rom[959] = 8'h0b ;
            rom[960] = 8'hf5 ;
            rom[961] = 8'h01 ;
            rom[962] = 8'h25 ;
            rom[963] = 8'h08 ;
            rom[964] = 8'h1d ;
            rom[965] = 8'h01 ;
            rom[966] = 8'hdd ;
            rom[967] = 8'h06 ;
            rom[968] = 8'hf4 ;
            rom[969] = 8'h03 ;
            rom[970] = 8'hfb ;
            rom[971] = 8'h1a ;
            rom[972] = 8'h0a ;
            rom[973] = 8'hfc ;
            rom[974] = 8'h1d ;
            rom[975] = 8'h05 ;
            rom[976] = 8'hfe ;
            rom[977] = 8'hb3 ;
            rom[978] = 8'h06 ;
            rom[979] = 8'hed ;
            rom[980] = 8'h07 ;
            rom[981] = 8'he0 ;
            rom[982] = 8'h02 ;
            rom[983] = 8'hfc ;
            rom[984] = 8'he6 ;
            rom[985] = 8'h0d ;
            rom[986] = 8'hf0 ;
            rom[987] = 8'h05 ;
            rom[988] = 8'hfd ;
            rom[989] = 8'hf8 ;
            rom[990] = 8'h16 ;
            rom[991] = 8'hfb ;
            rom[992] = 8'he6 ;
            rom[993] = 8'h00 ;
            rom[994] = 8'h24 ;
            rom[995] = 8'hff ;
            rom[996] = 8'hf3 ;
            rom[997] = 8'he4 ;
            rom[998] = 8'h14 ;
            rom[999] = 8'he9 ;
            rom[1000] = 8'hec ;
            rom[1001] = 8'hfe ;
            rom[1002] = 8'heb ;
            rom[1003] = 8'h02 ;
            rom[1004] = 8'hf8 ;
            rom[1005] = 8'h56 ;
            rom[1006] = 8'he7 ;
            rom[1007] = 8'h19 ;
            rom[1008] = 8'h03 ;
            rom[1009] = 8'hfa ;
            rom[1010] = 8'hf7 ;
            rom[1011] = 8'h14 ;
            rom[1012] = 8'hf2 ;
            rom[1013] = 8'he1 ;
            rom[1014] = 8'h27 ;
            rom[1015] = 8'h0f ;
            rom[1016] = 8'hfa ;
            rom[1017] = 8'hf0 ;
            rom[1018] = 8'hde ;
            rom[1019] = 8'h02 ;
            rom[1020] = 8'he3 ;
            rom[1021] = 8'h08 ;
            rom[1022] = 8'h07 ;
            rom[1023] = 8'h20 ;
            rom[1024] = 8'h0c ;
            rom[1025] = 8'hfc ;
            rom[1026] = 8'hdf ;
            rom[1027] = 8'h08 ;
            rom[1028] = 8'h00 ;
            rom[1029] = 8'h1c ;
            rom[1030] = 8'he5 ;
            rom[1031] = 8'h08 ;
            rom[1032] = 8'hec ;
            rom[1033] = 8'h0d ;
            rom[1034] = 8'h01 ;
            rom[1035] = 8'h0d ;
            rom[1036] = 8'h24 ;
            rom[1037] = 8'hdf ;
            rom[1038] = 8'h1d ;
            rom[1039] = 8'h0d ;
            rom[1040] = 8'hf5 ;
            rom[1041] = 8'hf5 ;
            rom[1042] = 8'hfe ;
            rom[1043] = 8'h11 ;
            rom[1044] = 8'h0f ;
            rom[1045] = 8'h39 ;
            rom[1046] = 8'h0c ;
            rom[1047] = 8'h00 ;
            rom[1048] = 8'hfa ;
            rom[1049] = 8'h0d ;
            rom[1050] = 8'he2 ;
            rom[1051] = 8'h02 ;
            rom[1052] = 8'hec ;
            rom[1053] = 8'h03 ;
            rom[1054] = 8'hfa ;
            rom[1055] = 8'he8 ;
            rom[1056] = 8'heb ;
            rom[1057] = 8'h0b ;
            rom[1058] = 8'h1c ;
            rom[1059] = 8'he7 ;
            rom[1060] = 8'he7 ;
            rom[1061] = 8'hfe ;
            rom[1062] = 8'hfb ;
            rom[1063] = 8'hfe ;
            rom[1064] = 8'h0b ;
            rom[1065] = 8'h15 ;
            rom[1066] = 8'hd2 ;
            rom[1067] = 8'hfd ;
            rom[1068] = 8'h00 ;
            rom[1069] = 8'h07 ;
            rom[1070] = 8'h0a ;
            rom[1071] = 8'hf6 ;
            rom[1072] = 8'h19 ;
            rom[1073] = 8'h0e ;
            rom[1074] = 8'hf7 ;
            rom[1075] = 8'h11 ;
            rom[1076] = 8'h16 ;
            rom[1077] = 8'hb6 ;
            rom[1078] = 8'hf1 ;
            rom[1079] = 8'h1a ;
            rom[1080] = 8'he2 ;
            rom[1081] = 8'h01 ;
            rom[1082] = 8'hf1 ;
            rom[1083] = 8'h17 ;
            rom[1084] = 8'he5 ;
            rom[1085] = 8'hcd ;
            rom[1086] = 8'h0b ;
            rom[1087] = 8'h35 ;
            rom[1088] = 8'h17 ;
            rom[1089] = 8'h05 ;
            rom[1090] = 8'hf8 ;
            rom[1091] = 8'h03 ;
            rom[1092] = 8'h00 ;
            rom[1093] = 8'h19 ;
            rom[1094] = 8'h03 ;
            rom[1095] = 8'h13 ;
            rom[1096] = 8'hee ;
            rom[1097] = 8'hf7 ;
            rom[1098] = 8'hf7 ;
            rom[1099] = 8'heb ;
            rom[1100] = 8'h28 ;
            rom[1101] = 8'h0f ;
            rom[1102] = 8'hfc ;
            rom[1103] = 8'hed ;
            rom[1104] = 8'hf5 ;
            rom[1105] = 8'h14 ;
            rom[1106] = 8'hbe ;
            rom[1107] = 8'h15 ;
            rom[1108] = 8'h09 ;
            rom[1109] = 8'h02 ;
            rom[1110] = 8'h1c ;
            rom[1111] = 8'h01 ;
            rom[1112] = 8'h02 ;
            rom[1113] = 8'h13 ;
            rom[1114] = 8'h08 ;
            rom[1115] = 8'hf4 ;
            rom[1116] = 8'h03 ;
            rom[1117] = 8'h0e ;
            rom[1118] = 8'h04 ;
            rom[1119] = 8'hef ;
            rom[1120] = 8'h0a ;
            rom[1121] = 8'hf0 ;
            rom[1122] = 8'hfe ;
            rom[1123] = 8'hff ;
            rom[1124] = 8'h07 ;
            rom[1125] = 8'h34 ;
            rom[1126] = 8'hf6 ;
            rom[1127] = 8'h10 ;
            rom[1128] = 8'h15 ;
            rom[1129] = 8'heb ;
            rom[1130] = 8'hf6 ;
            rom[1131] = 8'hff ;
            rom[1132] = 8'h07 ;
            rom[1133] = 8'hf3 ;
            rom[1134] = 8'h21 ;
            rom[1135] = 8'h0f ;
            rom[1136] = 8'h15 ;
            rom[1137] = 8'h14 ;
            rom[1138] = 8'h02 ;
            rom[1139] = 8'hcf ;
            rom[1140] = 8'h19 ;
            rom[1141] = 8'hf6 ;
            rom[1142] = 8'h18 ;
            rom[1143] = 8'h01 ;
            rom[1144] = 8'h19 ;
            rom[1145] = 8'heb ;
            rom[1146] = 8'hf8 ;
            rom[1147] = 8'hfb ;
            rom[1148] = 8'h05 ;
            rom[1149] = 8'h02 ;
            rom[1150] = 8'h20 ;
            rom[1151] = 8'h12 ;
            rom[1152] = 8'hd5 ;
            rom[1153] = 8'he1 ;
            rom[1154] = 8'hff ;
            rom[1155] = 8'h14 ;
            rom[1156] = 8'h1a ;
            rom[1157] = 8'h16 ;
            rom[1158] = 8'h02 ;
            rom[1159] = 8'he9 ;
            rom[1160] = 8'hf4 ;
            rom[1161] = 8'hfd ;
            rom[1162] = 8'hed ;
            rom[1163] = 8'h0a ;
            rom[1164] = 8'hfc ;
            rom[1165] = 8'hdd ;
            rom[1166] = 8'h02 ;
            rom[1167] = 8'hf7 ;
            rom[1168] = 8'hec ;
            rom[1169] = 8'hec ;
            rom[1170] = 8'hf6 ;
            rom[1171] = 8'h09 ;
            rom[1172] = 8'hf0 ;
            rom[1173] = 8'h01 ;
            rom[1174] = 8'h06 ;
            rom[1175] = 8'h20 ;
            rom[1176] = 8'hf7 ;
            rom[1177] = 8'h07 ;
            rom[1178] = 8'h03 ;
            rom[1179] = 8'h12 ;
            rom[1180] = 8'h07 ;
            rom[1181] = 8'hd4 ;
            rom[1182] = 8'h15 ;
            rom[1183] = 8'he3 ;
            rom[1184] = 8'h11 ;
            rom[1185] = 8'he3 ;
            rom[1186] = 8'hfc ;
            rom[1187] = 8'hfe ;
            rom[1188] = 8'h1d ;
            rom[1189] = 8'h16 ;
            rom[1190] = 8'hfd ;
            rom[1191] = 8'hec ;
            rom[1192] = 8'he3 ;
            rom[1193] = 8'h05 ;
            rom[1194] = 8'h12 ;
            rom[1195] = 8'h1a ;
            rom[1196] = 8'h0e ;
            rom[1197] = 8'h09 ;
            rom[1198] = 8'h02 ;
            rom[1199] = 8'hec ;
            rom[1200] = 8'hf7 ;
            rom[1201] = 8'h07 ;
            rom[1202] = 8'hfe ;
            rom[1203] = 8'hf0 ;
            rom[1204] = 8'hfe ;
            rom[1205] = 8'h06 ;
            rom[1206] = 8'h1e ;
            rom[1207] = 8'hfd ;
            rom[1208] = 8'h07 ;
            rom[1209] = 8'h08 ;
            rom[1210] = 8'h03 ;
            rom[1211] = 8'h11 ;
            rom[1212] = 8'hcd ;
            rom[1213] = 8'h03 ;
            rom[1214] = 8'h04 ;
            rom[1215] = 8'he7 ;
            rom[1216] = 8'hdf ;
            rom[1217] = 8'hec ;
            rom[1218] = 8'hff ;
            rom[1219] = 8'hf0 ;
            rom[1220] = 8'hf9 ;
            rom[1221] = 8'h01 ;
            rom[1222] = 8'h09 ;
            rom[1223] = 8'h0a ;
            rom[1224] = 8'h15 ;
            rom[1225] = 8'h21 ;
            rom[1226] = 8'he1 ;
            rom[1227] = 8'h10 ;
            rom[1228] = 8'hf0 ;
            rom[1229] = 8'heb ;
            rom[1230] = 8'hf2 ;
            rom[1231] = 8'h06 ;
            rom[1232] = 8'h05 ;
            rom[1233] = 8'h0d ;
            rom[1234] = 8'hf9 ;
            rom[1235] = 8'hed ;
            rom[1236] = 8'heb ;
            rom[1237] = 8'h0f ;
            rom[1238] = 8'hed ;
            rom[1239] = 8'hdc ;
            rom[1240] = 8'h04 ;
            rom[1241] = 8'h05 ;
            rom[1242] = 8'hff ;
            rom[1243] = 8'h23 ;
            rom[1244] = 8'hde ;
            rom[1245] = 8'h01 ;
            rom[1246] = 8'h06 ;
            rom[1247] = 8'h04 ;
            rom[1248] = 8'hfc ;
            rom[1249] = 8'h09 ;
            rom[1250] = 8'hfe ;
            rom[1251] = 8'h06 ;
            rom[1252] = 8'hdb ;
            rom[1253] = 8'hfe ;
            rom[1254] = 8'he2 ;
            rom[1255] = 8'h08 ;
            rom[1256] = 8'h2c ;
            rom[1257] = 8'h0a ;
            rom[1258] = 8'he7 ;
            rom[1259] = 8'hfc ;
            rom[1260] = 8'hed ;
            rom[1261] = 8'hfb ;
            rom[1262] = 8'hcf ;
            rom[1263] = 8'h19 ;
            rom[1264] = 8'h18 ;
            rom[1265] = 8'he1 ;
            rom[1266] = 8'h03 ;
            rom[1267] = 8'h01 ;
            rom[1268] = 8'h0e ;
            rom[1269] = 8'hfe ;
            rom[1270] = 8'hd0 ;
            rom[1271] = 8'h0f ;
            rom[1272] = 8'h14 ;
            rom[1273] = 8'hfa ;
            rom[1274] = 8'hf8 ;
            rom[1275] = 8'hf1 ;
            rom[1276] = 8'hfb ;
            rom[1277] = 8'h12 ;
            rom[1278] = 8'hfd ;
            rom[1279] = 8'hf9 ;
            rom[1280] = 8'h04 ;
            rom[1281] = 8'h0b ;
            rom[1282] = 8'h2c ;
            rom[1283] = 8'h05 ;
            rom[1284] = 8'h0a ;
            rom[1285] = 8'h2b ;
            rom[1286] = 8'h0b ;
            rom[1287] = 8'hee ;
            rom[1288] = 8'heb ;
            rom[1289] = 8'h12 ;
            rom[1290] = 8'hfe ;
            rom[1291] = 8'hf9 ;
            rom[1292] = 8'h08 ;
            rom[1293] = 8'hd0 ;
            rom[1294] = 8'h00 ;
            rom[1295] = 8'h1c ;
            rom[1296] = 8'he7 ;
            rom[1297] = 8'h0d ;
            rom[1298] = 8'hfc ;
            rom[1299] = 8'h19 ;
            rom[1300] = 8'h00 ;
            rom[1301] = 8'h09 ;
            rom[1302] = 8'h0b ;
            rom[1303] = 8'h15 ;
            rom[1304] = 8'hff ;
            rom[1305] = 8'hf6 ;
            rom[1306] = 8'hdc ;
            rom[1307] = 8'h01 ;
            rom[1308] = 8'h07 ;
            rom[1309] = 8'hf8 ;
            rom[1310] = 8'hcc ;
            rom[1311] = 8'he6 ;
            rom[1312] = 8'h13 ;
            rom[1313] = 8'hfb ;
            rom[1314] = 8'h04 ;
            rom[1315] = 8'h12 ;
            rom[1316] = 8'hfa ;
            rom[1317] = 8'hf6 ;
            rom[1318] = 8'h0d ;
            rom[1319] = 8'h11 ;
            rom[1320] = 8'h04 ;
            rom[1321] = 8'hef ;
            rom[1322] = 8'h02 ;
            rom[1323] = 8'h0e ;
            rom[1324] = 8'hf3 ;
            rom[1325] = 8'h18 ;
            rom[1326] = 8'h14 ;
            rom[1327] = 8'hf3 ;
            rom[1328] = 8'h16 ;
            rom[1329] = 8'h22 ;
            rom[1330] = 8'h0e ;
            rom[1331] = 8'hf5 ;
            rom[1332] = 8'h13 ;
            rom[1333] = 8'he8 ;
            rom[1334] = 8'he9 ;
            rom[1335] = 8'h11 ;
            rom[1336] = 8'h07 ;
            rom[1337] = 8'hc3 ;
            rom[1338] = 8'hea ;
            rom[1339] = 8'hff ;
            rom[1340] = 8'h21 ;
            rom[1341] = 8'he1 ;
            rom[1342] = 8'he5 ;
            rom[1343] = 8'h1f ;
            rom[1344] = 8'h04 ;
            rom[1345] = 8'h03 ;
            rom[1346] = 8'hfb ;
            rom[1347] = 8'h0f ;
            rom[1348] = 8'h03 ;
            rom[1349] = 8'hf3 ;
            rom[1350] = 8'h03 ;
            rom[1351] = 8'h0c ;
            rom[1352] = 8'h0e ;
            rom[1353] = 8'he0 ;
            rom[1354] = 8'h04 ;
            rom[1355] = 8'h07 ;
            rom[1356] = 8'h26 ;
            rom[1357] = 8'hd8 ;
            rom[1358] = 8'h24 ;
            rom[1359] = 8'h0a ;
            rom[1360] = 8'h15 ;
            rom[1361] = 8'h0c ;
            rom[1362] = 8'hf7 ;
            rom[1363] = 8'hfd ;
            rom[1364] = 8'h08 ;
            rom[1365] = 8'h13 ;
            rom[1366] = 8'hf1 ;
            rom[1367] = 8'hf5 ;
            rom[1368] = 8'h07 ;
            rom[1369] = 8'h14 ;
            rom[1370] = 8'heb ;
            rom[1371] = 8'h0a ;
            rom[1372] = 8'hea ;
            rom[1373] = 8'h21 ;
            rom[1374] = 8'h2d ;
            rom[1375] = 8'h0e ;
            rom[1376] = 8'he3 ;
            rom[1377] = 8'h0e ;
            rom[1378] = 8'hed ;
            rom[1379] = 8'hf8 ;
            rom[1380] = 8'h06 ;
            rom[1381] = 8'he2 ;
            rom[1382] = 8'h00 ;
            rom[1383] = 8'h02 ;
            rom[1384] = 8'hfd ;
            rom[1385] = 8'hf0 ;
            rom[1386] = 8'h0b ;
            rom[1387] = 8'hef ;
            rom[1388] = 8'hfb ;
            rom[1389] = 8'h17 ;
            rom[1390] = 8'h04 ;
            rom[1391] = 8'h04 ;
            rom[1392] = 8'h0f ;
            rom[1393] = 8'h06 ;
            rom[1394] = 8'h11 ;
            rom[1395] = 8'h05 ;
            rom[1396] = 8'h0e ;
            rom[1397] = 8'he9 ;
            rom[1398] = 8'h04 ;
            rom[1399] = 8'h00 ;
            rom[1400] = 8'hda ;
            rom[1401] = 8'hf3 ;
            rom[1402] = 8'h11 ;
            rom[1403] = 8'h23 ;
            rom[1404] = 8'he6 ;
            rom[1405] = 8'h0a ;
            rom[1406] = 8'h18 ;
            rom[1407] = 8'h00 ;
            rom[1408] = 8'h0e ;
            rom[1409] = 8'hfd ;
            rom[1410] = 8'hdc ;
            rom[1411] = 8'hf8 ;
            rom[1412] = 8'h03 ;
            rom[1413] = 8'heb ;
            rom[1414] = 8'hf6 ;
            rom[1415] = 8'hfe ;
            rom[1416] = 8'h05 ;
            rom[1417] = 8'hfc ;
            rom[1418] = 8'h06 ;
            rom[1419] = 8'h1d ;
            rom[1420] = 8'h07 ;
            rom[1421] = 8'hff ;
            rom[1422] = 8'he0 ;
            rom[1423] = 8'hfe ;
            rom[1424] = 8'h07 ;
            rom[1425] = 8'h04 ;
            rom[1426] = 8'h0e ;
            rom[1427] = 8'hf0 ;
            rom[1428] = 8'h17 ;
            rom[1429] = 8'h07 ;
            rom[1430] = 8'he4 ;
            rom[1431] = 8'h13 ;
            rom[1432] = 8'hff ;
            rom[1433] = 8'hf7 ;
            rom[1434] = 8'hed ;
            rom[1435] = 8'h0e ;
            rom[1436] = 8'h0b ;
            rom[1437] = 8'h0e ;
            rom[1438] = 8'h02 ;
            rom[1439] = 8'h18 ;
            rom[1440] = 8'h07 ;
            rom[1441] = 8'h0a ;
            rom[1442] = 8'hcb ;
            rom[1443] = 8'hfb ;
            rom[1444] = 8'h0a ;
            rom[1445] = 8'hea ;
            rom[1446] = 8'he1 ;
            rom[1447] = 8'h10 ;
            rom[1448] = 8'hf9 ;
            rom[1449] = 8'h11 ;
            rom[1450] = 8'hf0 ;
            rom[1451] = 8'h0f ;
            rom[1452] = 8'hf1 ;
            rom[1453] = 8'h02 ;
            rom[1454] = 8'h03 ;
            rom[1455] = 8'h11 ;
            rom[1456] = 8'hfc ;
            rom[1457] = 8'hd2 ;
            rom[1458] = 8'hf2 ;
            rom[1459] = 8'hef ;
            rom[1460] = 8'hdb ;
            rom[1461] = 8'h12 ;
            rom[1462] = 8'hf3 ;
            rom[1463] = 8'hf9 ;
            rom[1464] = 8'hea ;
            rom[1465] = 8'h12 ;
            rom[1466] = 8'h04 ;
            rom[1467] = 8'h14 ;
            rom[1468] = 8'hfc ;
            rom[1469] = 8'hfb ;
            rom[1470] = 8'h13 ;
            rom[1471] = 8'h01 ;
            rom[1472] = 8'hf2 ;
            rom[1473] = 8'hf7 ;
            rom[1474] = 8'hc1 ;
            rom[1475] = 8'h0d ;
            rom[1476] = 8'h14 ;
            rom[1477] = 8'h02 ;
            rom[1478] = 8'h1d ;
            rom[1479] = 8'h1d ;
            rom[1480] = 8'hf6 ;
            rom[1481] = 8'hfd ;
            rom[1482] = 8'he7 ;
            rom[1483] = 8'hf5 ;
            rom[1484] = 8'hf8 ;
            rom[1485] = 8'h03 ;
            rom[1486] = 8'h25 ;
            rom[1487] = 8'hec ;
            rom[1488] = 8'h14 ;
            rom[1489] = 8'h09 ;
            rom[1490] = 8'hf7 ;
            rom[1491] = 8'h14 ;
            rom[1492] = 8'h19 ;
            rom[1493] = 8'h06 ;
            rom[1494] = 8'h0b ;
            rom[1495] = 8'h19 ;
            rom[1496] = 8'h09 ;
            rom[1497] = 8'h16 ;
            rom[1498] = 8'hf7 ;
            rom[1499] = 8'h18 ;
            rom[1500] = 8'hed ;
            rom[1501] = 8'h2a ;
            rom[1502] = 8'h21 ;
            rom[1503] = 8'hf4 ;
            rom[1504] = 8'hea ;
            rom[1505] = 8'hfc ;
            rom[1506] = 8'he2 ;
            rom[1507] = 8'h11 ;
            rom[1508] = 8'hf7 ;
            rom[1509] = 8'he5 ;
            rom[1510] = 8'hfc ;
            rom[1511] = 8'h0f ;
            rom[1512] = 8'h0f ;
            rom[1513] = 8'h01 ;
            rom[1514] = 8'h01 ;
            rom[1515] = 8'h09 ;
            rom[1516] = 8'hfc ;
            rom[1517] = 8'h22 ;
            rom[1518] = 8'hf6 ;
            rom[1519] = 8'h0f ;
            rom[1520] = 8'hfa ;
            rom[1521] = 8'h07 ;
            rom[1522] = 8'h12 ;
            rom[1523] = 8'hf6 ;
            rom[1524] = 8'h02 ;
            rom[1525] = 8'hdd ;
            rom[1526] = 8'h11 ;
            rom[1527] = 8'h03 ;
            rom[1528] = 8'he3 ;
            rom[1529] = 8'hea ;
            rom[1530] = 8'h16 ;
            rom[1531] = 8'h2f ;
            rom[1532] = 8'hd0 ;
            rom[1533] = 8'hf8 ;
            rom[1534] = 8'hf9 ;
            rom[1535] = 8'h0d ;
            rom[1536] = 8'hf3 ;
            rom[1537] = 8'hce ;
            rom[1538] = 8'h11 ;
            rom[1539] = 8'hfd ;
            rom[1540] = 8'h02 ;
            rom[1541] = 8'h04 ;
            rom[1542] = 8'hf6 ;
            rom[1543] = 8'hf5 ;
            rom[1544] = 8'hc6 ;
            rom[1545] = 8'h0f ;
            rom[1546] = 8'hfa ;
            rom[1547] = 8'h04 ;
            rom[1548] = 8'h03 ;
            rom[1549] = 8'hf2 ;
            rom[1550] = 8'hde ;
            rom[1551] = 8'h06 ;
            rom[1552] = 8'h07 ;
            rom[1553] = 8'hf3 ;
            rom[1554] = 8'he1 ;
            rom[1555] = 8'h0c ;
            rom[1556] = 8'h07 ;
            rom[1557] = 8'hfa ;
            rom[1558] = 8'h11 ;
            rom[1559] = 8'hfa ;
            rom[1560] = 8'h1d ;
            rom[1561] = 8'h09 ;
            rom[1562] = 8'hef ;
            rom[1563] = 8'h00 ;
            rom[1564] = 8'h07 ;
            rom[1565] = 8'hef ;
            rom[1566] = 8'hef ;
            rom[1567] = 8'he3 ;
            rom[1568] = 8'h0e ;
            rom[1569] = 8'he8 ;
            rom[1570] = 8'hdf ;
            rom[1571] = 8'h16 ;
            rom[1572] = 8'hfd ;
            rom[1573] = 8'h03 ;
            rom[1574] = 8'hf3 ;
            rom[1575] = 8'h06 ;
            rom[1576] = 8'hfa ;
            rom[1577] = 8'he0 ;
            rom[1578] = 8'hee ;
            rom[1579] = 8'h00 ;
            rom[1580] = 8'he7 ;
            rom[1581] = 8'hfe ;
            rom[1582] = 8'h1f ;
            rom[1583] = 8'h27 ;
            rom[1584] = 8'h0b ;
            rom[1585] = 8'h20 ;
            rom[1586] = 8'h0e ;
            rom[1587] = 8'hde ;
            rom[1588] = 8'hf5 ;
            rom[1589] = 8'hea ;
            rom[1590] = 8'h0c ;
            rom[1591] = 8'h05 ;
            rom[1592] = 8'he8 ;
            rom[1593] = 8'hec ;
            rom[1594] = 8'hd1 ;
            rom[1595] = 8'hfb ;
            rom[1596] = 8'h01 ;
            rom[1597] = 8'hee ;
            rom[1598] = 8'h0e ;
            rom[1599] = 8'hec ;
            rom[1600] = 8'hef ;
            rom[1601] = 8'h08 ;
            rom[1602] = 8'hfd ;
            rom[1603] = 8'h00 ;
            rom[1604] = 8'h10 ;
            rom[1605] = 8'hf9 ;
            rom[1606] = 8'h08 ;
            rom[1607] = 8'h18 ;
            rom[1608] = 8'hff ;
            rom[1609] = 8'h22 ;
            rom[1610] = 8'hae ;
            rom[1611] = 8'h02 ;
            rom[1612] = 8'he1 ;
            rom[1613] = 8'hea ;
            rom[1614] = 8'h05 ;
            rom[1615] = 8'h00 ;
            rom[1616] = 8'h1e ;
            rom[1617] = 8'h0d ;
            rom[1618] = 8'hf6 ;
            rom[1619] = 8'he5 ;
            rom[1620] = 8'h03 ;
            rom[1621] = 8'h0e ;
            rom[1622] = 8'hfc ;
            rom[1623] = 8'hfa ;
            rom[1624] = 8'h0c ;
            rom[1625] = 8'h0e ;
            rom[1626] = 8'h1e ;
            rom[1627] = 8'hff ;
            rom[1628] = 8'he6 ;
            rom[1629] = 8'h2a ;
            rom[1630] = 8'h03 ;
            rom[1631] = 8'he3 ;
            rom[1632] = 8'h05 ;
            rom[1633] = 8'hf8 ;
            rom[1634] = 8'hff ;
            rom[1635] = 8'h02 ;
            rom[1636] = 8'hd7 ;
            rom[1637] = 8'h05 ;
            rom[1638] = 8'he3 ;
            rom[1639] = 8'h14 ;
            rom[1640] = 8'h20 ;
            rom[1641] = 8'hd3 ;
            rom[1642] = 8'he7 ;
            rom[1643] = 8'hf4 ;
            rom[1644] = 8'hf1 ;
            rom[1645] = 8'h16 ;
            rom[1646] = 8'hd8 ;
            rom[1647] = 8'h07 ;
            rom[1648] = 8'h07 ;
            rom[1649] = 8'he9 ;
            rom[1650] = 8'hed ;
            rom[1651] = 8'h06 ;
            rom[1652] = 8'hf5 ;
            rom[1653] = 8'h00 ;
            rom[1654] = 8'he5 ;
            rom[1655] = 8'h01 ;
            rom[1656] = 8'h02 ;
            rom[1657] = 8'h0a ;
            rom[1658] = 8'hfc ;
            rom[1659] = 8'h0f ;
            rom[1660] = 8'h0e ;
            rom[1661] = 8'h11 ;
            rom[1662] = 8'hfd ;
            rom[1663] = 8'h00 ;
            rom[1664] = 8'h00 ;
            rom[1665] = 8'h16 ;
            rom[1666] = 8'h0a ;
            rom[1667] = 8'hf4 ;
            rom[1668] = 8'h06 ;
            rom[1669] = 8'he4 ;
            rom[1670] = 8'h17 ;
            rom[1671] = 8'h0a ;
            rom[1672] = 8'h03 ;
            rom[1673] = 8'hed ;
            rom[1674] = 8'hde ;
            rom[1675] = 8'hf2 ;
            rom[1676] = 8'h0e ;
            rom[1677] = 8'h09 ;
            rom[1678] = 8'h0a ;
            rom[1679] = 8'h1a ;
            rom[1680] = 8'h18 ;
            rom[1681] = 8'h17 ;
            rom[1682] = 8'h0c ;
            rom[1683] = 8'he3 ;
            rom[1684] = 8'h0c ;
            rom[1685] = 8'hfa ;
            rom[1686] = 8'h04 ;
            rom[1687] = 8'hfe ;
            rom[1688] = 8'hf2 ;
            rom[1689] = 8'hf9 ;
            rom[1690] = 8'h12 ;
            rom[1691] = 8'h0a ;
            rom[1692] = 8'hed ;
            rom[1693] = 8'hee ;
            rom[1694] = 8'hf2 ;
            rom[1695] = 8'h01 ;
            rom[1696] = 8'hf1 ;
            rom[1697] = 8'h12 ;
            rom[1698] = 8'hd3 ;
            rom[1699] = 8'hf0 ;
            rom[1700] = 8'h00 ;
            rom[1701] = 8'he7 ;
            rom[1702] = 8'hda ;
            rom[1703] = 8'he9 ;
            rom[1704] = 8'hf8 ;
            rom[1705] = 8'hb1 ;
            rom[1706] = 8'h1b ;
            rom[1707] = 8'he0 ;
            rom[1708] = 8'h0a ;
            rom[1709] = 8'hfb ;
            rom[1710] = 8'hc9 ;
            rom[1711] = 8'h0a ;
            rom[1712] = 8'h06 ;
            rom[1713] = 8'hf3 ;
            rom[1714] = 8'h00 ;
            rom[1715] = 8'he6 ;
            rom[1716] = 8'h12 ;
            rom[1717] = 8'h0e ;
            rom[1718] = 8'h1a ;
            rom[1719] = 8'h13 ;
            rom[1720] = 8'he6 ;
            rom[1721] = 8'h05 ;
            rom[1722] = 8'hfa ;
            rom[1723] = 8'h1f ;
            rom[1724] = 8'h02 ;
            rom[1725] = 8'h12 ;
            rom[1726] = 8'h1a ;
            rom[1727] = 8'h0f ;
            rom[1728] = 8'hef ;
            rom[1729] = 8'h20 ;
            rom[1730] = 8'hcb ;
            rom[1731] = 8'hf8 ;
            rom[1732] = 8'hfd ;
            rom[1733] = 8'he1 ;
            rom[1734] = 8'h11 ;
            rom[1735] = 8'h0a ;
            rom[1736] = 8'h01 ;
            rom[1737] = 8'hf6 ;
            rom[1738] = 8'hda ;
            rom[1739] = 8'hf5 ;
            rom[1740] = 8'hff ;
            rom[1741] = 8'he5 ;
            rom[1742] = 8'hfd ;
            rom[1743] = 8'hfc ;
            rom[1744] = 8'hfe ;
            rom[1745] = 8'h11 ;
            rom[1746] = 8'he6 ;
            rom[1747] = 8'hff ;
            rom[1748] = 8'h17 ;
            rom[1749] = 8'h06 ;
            rom[1750] = 8'h00 ;
            rom[1751] = 8'hf2 ;
            rom[1752] = 8'he9 ;
            rom[1753] = 8'h35 ;
            rom[1754] = 8'he7 ;
            rom[1755] = 8'h13 ;
            rom[1756] = 8'hea ;
            rom[1757] = 8'h06 ;
            rom[1758] = 8'h18 ;
            rom[1759] = 8'hf2 ;
            rom[1760] = 8'hef ;
            rom[1761] = 8'hff ;
            rom[1762] = 8'hbd ;
            rom[1763] = 8'hf2 ;
            rom[1764] = 8'hf1 ;
            rom[1765] = 8'hea ;
            rom[1766] = 8'hee ;
            rom[1767] = 8'h0c ;
            rom[1768] = 8'h24 ;
            rom[1769] = 8'hf6 ;
            rom[1770] = 8'h21 ;
            rom[1771] = 8'hdc ;
            rom[1772] = 8'hf4 ;
            rom[1773] = 8'h13 ;
            rom[1774] = 8'h09 ;
            rom[1775] = 8'h06 ;
            rom[1776] = 8'h09 ;
            rom[1777] = 8'hfc ;
            rom[1778] = 8'h17 ;
            rom[1779] = 8'hd5 ;
            rom[1780] = 8'hf6 ;
            rom[1781] = 8'hfc ;
            rom[1782] = 8'he0 ;
            rom[1783] = 8'h07 ;
            rom[1784] = 8'he2 ;
            rom[1785] = 8'hee ;
            rom[1786] = 8'h06 ;
            rom[1787] = 8'h13 ;
            rom[1788] = 8'hf4 ;
            rom[1789] = 8'heb ;
            rom[1790] = 8'hf7 ;
            rom[1791] = 8'h0f ;
            rom[1792] = 8'h14 ;
            rom[1793] = 8'h04 ;
            rom[1794] = 8'hf0 ;
            rom[1795] = 8'h1c ;
            rom[1796] = 8'he9 ;
            rom[1797] = 8'h02 ;
            rom[1798] = 8'hfb ;
            rom[1799] = 8'h0b ;
            rom[1800] = 8'he7 ;
            rom[1801] = 8'hd7 ;
            rom[1802] = 8'h08 ;
            rom[1803] = 8'h00 ;
            rom[1804] = 8'hfb ;
            rom[1805] = 8'hd3 ;
            rom[1806] = 8'hee ;
            rom[1807] = 8'h00 ;
            rom[1808] = 8'h0e ;
            rom[1809] = 8'h17 ;
            rom[1810] = 8'h00 ;
            rom[1811] = 8'hfb ;
            rom[1812] = 8'h08 ;
            rom[1813] = 8'h22 ;
            rom[1814] = 8'hf5 ;
            rom[1815] = 8'h0b ;
            rom[1816] = 8'hff ;
            rom[1817] = 8'h10 ;
            rom[1818] = 8'hf8 ;
            rom[1819] = 8'h19 ;
            rom[1820] = 8'he2 ;
            rom[1821] = 8'h19 ;
            rom[1822] = 8'hff ;
            rom[1823] = 8'hfa ;
            rom[1824] = 8'hc6 ;
            rom[1825] = 8'hf2 ;
            rom[1826] = 8'hf1 ;
            rom[1827] = 8'hf9 ;
            rom[1828] = 8'hfe ;
            rom[1829] = 8'hbe ;
            rom[1830] = 8'h0c ;
            rom[1831] = 8'hfb ;
            rom[1832] = 8'hea ;
            rom[1833] = 8'hf8 ;
            rom[1834] = 8'hdc ;
            rom[1835] = 8'h10 ;
            rom[1836] = 8'hf3 ;
            rom[1837] = 8'h1f ;
            rom[1838] = 8'h16 ;
            rom[1839] = 8'hd7 ;
            rom[1840] = 8'h1a ;
            rom[1841] = 8'hed ;
            rom[1842] = 8'h09 ;
            rom[1843] = 8'hd9 ;
            rom[1844] = 8'hf6 ;
            rom[1845] = 8'hef ;
            rom[1846] = 8'hee ;
            rom[1847] = 8'h0b ;
            rom[1848] = 8'hf2 ;
            rom[1849] = 8'hf5 ;
            rom[1850] = 8'hf7 ;
            rom[1851] = 8'h0d ;
            rom[1852] = 8'hf2 ;
            rom[1853] = 8'he3 ;
            rom[1854] = 8'he5 ;
            rom[1855] = 8'h1b ;
            rom[1856] = 8'h15 ;
            rom[1857] = 8'h1a ;
            rom[1858] = 8'h1d ;
            rom[1859] = 8'he3 ;
            rom[1860] = 8'h16 ;
            rom[1861] = 8'h13 ;
            rom[1862] = 8'hee ;
            rom[1863] = 8'hf9 ;
            rom[1864] = 8'h10 ;
            rom[1865] = 8'h09 ;
            rom[1866] = 8'hfa ;
            rom[1867] = 8'he6 ;
            rom[1868] = 8'h09 ;
            rom[1869] = 8'hce ;
            rom[1870] = 8'h11 ;
            rom[1871] = 8'he2 ;
            rom[1872] = 8'hef ;
            rom[1873] = 8'h09 ;
            rom[1874] = 8'he2 ;
            rom[1875] = 8'h01 ;
            rom[1876] = 8'he8 ;
            rom[1877] = 8'hdd ;
            rom[1878] = 8'h02 ;
            rom[1879] = 8'hf4 ;
            rom[1880] = 8'h03 ;
            rom[1881] = 8'h0f ;
            rom[1882] = 8'h07 ;
            rom[1883] = 8'h06 ;
            rom[1884] = 8'h08 ;
            rom[1885] = 8'h17 ;
            rom[1886] = 8'he8 ;
            rom[1887] = 8'h0e ;
            rom[1888] = 8'hfa ;
            rom[1889] = 8'hf2 ;
            rom[1890] = 8'hf5 ;
            rom[1891] = 8'h1c ;
            rom[1892] = 8'hea ;
            rom[1893] = 8'hf5 ;
            rom[1894] = 8'hf4 ;
            rom[1895] = 8'hfa ;
            rom[1896] = 8'h0d ;
            rom[1897] = 8'hd8 ;
            rom[1898] = 8'h16 ;
            rom[1899] = 8'h0f ;
            rom[1900] = 8'hc1 ;
            rom[1901] = 8'h0f ;
            rom[1902] = 8'h04 ;
            rom[1903] = 8'hb9 ;
            rom[1904] = 8'h2b ;
            rom[1905] = 8'h1d ;
            rom[1906] = 8'he3 ;
            rom[1907] = 8'hea ;
            rom[1908] = 8'hf7 ;
            rom[1909] = 8'h10 ;
            rom[1910] = 8'hf1 ;
            rom[1911] = 8'h11 ;
            rom[1912] = 8'h0a ;
            rom[1913] = 8'hf6 ;
            rom[1914] = 8'he4 ;
            rom[1915] = 8'hed ;
            rom[1916] = 8'h03 ;
            rom[1917] = 8'hff ;
            rom[1918] = 8'hff ;
            rom[1919] = 8'hfe ;
            rom[1920] = 8'he4 ;
            rom[1921] = 8'he3 ;
            rom[1922] = 8'h0f ;
            rom[1923] = 8'h05 ;
            rom[1924] = 8'h20 ;
            rom[1925] = 8'h12 ;
            rom[1926] = 8'hf3 ;
            rom[1927] = 8'hf0 ;
            rom[1928] = 8'hc7 ;
            rom[1929] = 8'h06 ;
            rom[1930] = 8'h02 ;
            rom[1931] = 8'h28 ;
            rom[1932] = 8'h02 ;
            rom[1933] = 8'hfe ;
            rom[1934] = 8'h06 ;
            rom[1935] = 8'h01 ;
            rom[1936] = 8'hed ;
            rom[1937] = 8'h09 ;
            rom[1938] = 8'h2e ;
            rom[1939] = 8'h04 ;
            rom[1940] = 8'h18 ;
            rom[1941] = 8'hd5 ;
            rom[1942] = 8'hf6 ;
            rom[1943] = 8'h1b ;
            rom[1944] = 8'hde ;
            rom[1945] = 8'hd8 ;
            rom[1946] = 8'hfa ;
            rom[1947] = 8'h0d ;
            rom[1948] = 8'h0a ;
            rom[1949] = 8'h0a ;
            rom[1950] = 8'hfc ;
            rom[1951] = 8'h17 ;
            rom[1952] = 8'he4 ;
            rom[1953] = 8'hec ;
            rom[1954] = 8'h05 ;
            rom[1955] = 8'hd9 ;
            rom[1956] = 8'h28 ;
            rom[1957] = 8'hf8 ;
            rom[1958] = 8'h20 ;
            rom[1959] = 8'h0d ;
            rom[1960] = 8'h18 ;
            rom[1961] = 8'hff ;
            rom[1962] = 8'hf5 ;
            rom[1963] = 8'h0b ;
            rom[1964] = 8'h00 ;
            rom[1965] = 8'h2f ;
            rom[1966] = 8'he7 ;
            rom[1967] = 8'h10 ;
            rom[1968] = 8'h16 ;
            rom[1969] = 8'he2 ;
            rom[1970] = 8'hea ;
            rom[1971] = 8'h06 ;
            rom[1972] = 8'hee ;
            rom[1973] = 8'hf0 ;
            rom[1974] = 8'h1f ;
            rom[1975] = 8'hfa ;
            rom[1976] = 8'h06 ;
            rom[1977] = 8'h07 ;
            rom[1978] = 8'hcd ;
            rom[1979] = 8'h16 ;
            rom[1980] = 8'hfd ;
            rom[1981] = 8'hfd ;
            rom[1982] = 8'h16 ;
            rom[1983] = 8'hfd ;
            rom[1984] = 8'h22 ;
            rom[1985] = 8'h05 ;
            rom[1986] = 8'hfd ;
            rom[1987] = 8'h15 ;
            rom[1988] = 8'h14 ;
            rom[1989] = 8'hfb ;
            rom[1990] = 8'h01 ;
            rom[1991] = 8'h08 ;
            rom[1992] = 8'hfd ;
            rom[1993] = 8'hf3 ;
            rom[1994] = 8'h0b ;
            rom[1995] = 8'hf9 ;
            rom[1996] = 8'hf2 ;
            rom[1997] = 8'hfd ;
            rom[1998] = 8'h0f ;
            rom[1999] = 8'h00 ;
            rom[2000] = 8'hff ;
            rom[2001] = 8'hfd ;
            rom[2002] = 8'hb7 ;
            rom[2003] = 8'hd7 ;
            rom[2004] = 8'h00 ;
            rom[2005] = 8'hf1 ;
            rom[2006] = 8'h0c ;
            rom[2007] = 8'hde ;
            rom[2008] = 8'hed ;
            rom[2009] = 8'h0b ;
            rom[2010] = 8'h22 ;
            rom[2011] = 8'h0c ;
            rom[2012] = 8'h1b ;
            rom[2013] = 8'h1a ;
            rom[2014] = 8'hf0 ;
            rom[2015] = 8'hff ;
            rom[2016] = 8'h10 ;
            rom[2017] = 8'hd6 ;
            rom[2018] = 8'h08 ;
            rom[2019] = 8'h00 ;
            rom[2020] = 8'hf0 ;
            rom[2021] = 8'hf9 ;
            rom[2022] = 8'hfc ;
            rom[2023] = 8'hd8 ;
            rom[2024] = 8'he9 ;
            rom[2025] = 8'hf1 ;
            rom[2026] = 8'h31 ;
            rom[2027] = 8'hfe ;
            rom[2028] = 8'hf5 ;
            rom[2029] = 8'h0b ;
            rom[2030] = 8'h10 ;
            rom[2031] = 8'h08 ;
            rom[2032] = 8'h0e ;
            rom[2033] = 8'hf3 ;
            rom[2034] = 8'hf1 ;
            rom[2035] = 8'h04 ;
            rom[2036] = 8'hed ;
            rom[2037] = 8'h0e ;
            rom[2038] = 8'h16 ;
            rom[2039] = 8'h14 ;
            rom[2040] = 8'heb ;
            rom[2041] = 8'h2b ;
            rom[2042] = 8'h0a ;
            rom[2043] = 8'hdf ;
            rom[2044] = 8'hf9 ;
            rom[2045] = 8'h0a ;
            rom[2046] = 8'h0f ;
            rom[2047] = 8'hf1 ;
            rom[2048] = 8'h18 ;
            rom[2049] = 8'h0a ;
            rom[2050] = 8'hf4 ;
            rom[2051] = 8'h0d ;
            rom[2052] = 8'he6 ;
            rom[2053] = 8'h1c ;
            rom[2054] = 8'hde ;
            rom[2055] = 8'hbd ;
            rom[2056] = 8'hf0 ;
            rom[2057] = 8'h07 ;
            rom[2058] = 8'hf5 ;
            rom[2059] = 8'h03 ;
            rom[2060] = 8'hcf ;
            rom[2061] = 8'he9 ;
            rom[2062] = 8'h33 ;
            rom[2063] = 8'hf4 ;
            rom[2064] = 8'heb ;
            rom[2065] = 8'hff ;
            rom[2066] = 8'he8 ;
            rom[2067] = 8'he4 ;
            rom[2068] = 8'h0f ;
            rom[2069] = 8'hf2 ;
            rom[2070] = 8'h0f ;
            rom[2071] = 8'hfe ;
            rom[2072] = 8'hf9 ;
            rom[2073] = 8'h01 ;
            rom[2074] = 8'h0a ;
            rom[2075] = 8'hee ;
            rom[2076] = 8'hf9 ;
            rom[2077] = 8'h06 ;
            rom[2078] = 8'hfc ;
            rom[2079] = 8'hf3 ;
            rom[2080] = 8'h09 ;
            rom[2081] = 8'he9 ;
            rom[2082] = 8'hfb ;
            rom[2083] = 8'h00 ;
            rom[2084] = 8'he9 ;
            rom[2085] = 8'h04 ;
            rom[2086] = 8'h14 ;
            rom[2087] = 8'hf3 ;
            rom[2088] = 8'hfd ;
            rom[2089] = 8'hdd ;
            rom[2090] = 8'he7 ;
            rom[2091] = 8'h16 ;
            rom[2092] = 8'h06 ;
            rom[2093] = 8'hed ;
            rom[2094] = 8'hf5 ;
            rom[2095] = 8'hee ;
            rom[2096] = 8'h01 ;
            rom[2097] = 8'h2b ;
            rom[2098] = 8'hfb ;
            rom[2099] = 8'hfc ;
            rom[2100] = 8'hee ;
            rom[2101] = 8'he7 ;
            rom[2102] = 8'hed ;
            rom[2103] = 8'hcb ;
            rom[2104] = 8'h15 ;
            rom[2105] = 8'h18 ;
            rom[2106] = 8'he7 ;
            rom[2107] = 8'he1 ;
            rom[2108] = 8'hfd ;
            rom[2109] = 8'h0f ;
            rom[2110] = 8'h0c ;
            rom[2111] = 8'hce ;
            rom[2112] = 8'h11 ;
            rom[2113] = 8'he9 ;
            rom[2114] = 8'hf0 ;
            rom[2115] = 8'hc9 ;
            rom[2116] = 8'h0b ;
            rom[2117] = 8'hfb ;
            rom[2118] = 8'hdd ;
            rom[2119] = 8'he7 ;
            rom[2120] = 8'h02 ;
            rom[2121] = 8'hf2 ;
            rom[2122] = 8'hf1 ;
            rom[2123] = 8'hf9 ;
            rom[2124] = 8'h0d ;
            rom[2125] = 8'he4 ;
            rom[2126] = 8'hef ;
            rom[2127] = 8'h05 ;
            rom[2128] = 8'hfa ;
            rom[2129] = 8'h0c ;
            rom[2130] = 8'hfc ;
            rom[2131] = 8'h02 ;
            rom[2132] = 8'h04 ;
            rom[2133] = 8'hf2 ;
            rom[2134] = 8'h15 ;
            rom[2135] = 8'h09 ;
            rom[2136] = 8'hf6 ;
            rom[2137] = 8'hf1 ;
            rom[2138] = 8'hdf ;
            rom[2139] = 8'hed ;
            rom[2140] = 8'h06 ;
            rom[2141] = 8'hfe ;
            rom[2142] = 8'hf1 ;
            rom[2143] = 8'he8 ;
            rom[2144] = 8'h16 ;
            rom[2145] = 8'hfb ;
            rom[2146] = 8'hf3 ;
            rom[2147] = 8'h10 ;
            rom[2148] = 8'h1e ;
            rom[2149] = 8'h0e ;
            rom[2150] = 8'hfc ;
            rom[2151] = 8'hee ;
            rom[2152] = 8'h1a ;
            rom[2153] = 8'hdd ;
            rom[2154] = 8'hf4 ;
            rom[2155] = 8'h07 ;
            rom[2156] = 8'hfc ;
            rom[2157] = 8'h10 ;
            rom[2158] = 8'h0f ;
            rom[2159] = 8'hfe ;
            rom[2160] = 8'hf7 ;
            rom[2161] = 8'hf6 ;
            rom[2162] = 8'hf6 ;
            rom[2163] = 8'h16 ;
            rom[2164] = 8'hf3 ;
            rom[2165] = 8'hfb ;
            rom[2166] = 8'he6 ;
            rom[2167] = 8'hf3 ;
            rom[2168] = 8'h07 ;
            rom[2169] = 8'hf8 ;
            rom[2170] = 8'hc6 ;
            rom[2171] = 8'h15 ;
            rom[2172] = 8'h0c ;
            rom[2173] = 8'hee ;
            rom[2174] = 8'h1b ;
            rom[2175] = 8'hf2 ;
            rom[2176] = 8'h10 ;
            rom[2177] = 8'he2 ;
            rom[2178] = 8'hfe ;
            rom[2179] = 8'h01 ;
            rom[2180] = 8'h0b ;
            rom[2181] = 8'he3 ;
            rom[2182] = 8'hd8 ;
            rom[2183] = 8'h05 ;
            rom[2184] = 8'h0c ;
            rom[2185] = 8'hf3 ;
            rom[2186] = 8'hfc ;
            rom[2187] = 8'h0b ;
            rom[2188] = 8'h13 ;
            rom[2189] = 8'hfb ;
            rom[2190] = 8'hfa ;
            rom[2191] = 8'h12 ;
            rom[2192] = 8'h05 ;
            rom[2193] = 8'h05 ;
            rom[2194] = 8'hd3 ;
            rom[2195] = 8'h14 ;
            rom[2196] = 8'hfd ;
            rom[2197] = 8'hd8 ;
            rom[2198] = 8'h17 ;
            rom[2199] = 8'hf4 ;
            rom[2200] = 8'h05 ;
            rom[2201] = 8'hfe ;
            rom[2202] = 8'h08 ;
            rom[2203] = 8'h0b ;
            rom[2204] = 8'h0f ;
            rom[2205] = 8'hf1 ;
            rom[2206] = 8'hf9 ;
            rom[2207] = 8'hdc ;
            rom[2208] = 8'hf0 ;
            rom[2209] = 8'hf8 ;
            rom[2210] = 8'h0c ;
            rom[2211] = 8'h03 ;
            rom[2212] = 8'he5 ;
            rom[2213] = 8'he6 ;
            rom[2214] = 8'hf5 ;
            rom[2215] = 8'hf7 ;
            rom[2216] = 8'hf9 ;
            rom[2217] = 8'hf8 ;
            rom[2218] = 8'h14 ;
            rom[2219] = 8'hfd ;
            rom[2220] = 8'heb ;
            rom[2221] = 8'h15 ;
            rom[2222] = 8'hf3 ;
            rom[2223] = 8'h17 ;
            rom[2224] = 8'hf6 ;
            rom[2225] = 8'h05 ;
            rom[2226] = 8'h10 ;
            rom[2227] = 8'hff ;
            rom[2228] = 8'hfe ;
            rom[2229] = 8'hd4 ;
            rom[2230] = 8'h06 ;
            rom[2231] = 8'h16 ;
            rom[2232] = 8'he9 ;
            rom[2233] = 8'hfb ;
            rom[2234] = 8'hf1 ;
            rom[2235] = 8'h02 ;
            rom[2236] = 8'hdf ;
            rom[2237] = 8'hf3 ;
            rom[2238] = 8'h10 ;
            rom[2239] = 8'hdc ;
            rom[2240] = 8'h1d ;
            rom[2241] = 8'he0 ;
            rom[2242] = 8'hf0 ;
            rom[2243] = 8'h07 ;
            rom[2244] = 8'h07 ;
            rom[2245] = 8'h15 ;
            rom[2246] = 8'hc7 ;
            rom[2247] = 8'hf1 ;
            rom[2248] = 8'h00 ;
            rom[2249] = 8'hf4 ;
            rom[2250] = 8'h02 ;
            rom[2251] = 8'h04 ;
            rom[2252] = 8'h1a ;
            rom[2253] = 8'he1 ;
            rom[2254] = 8'h26 ;
            rom[2255] = 8'hfe ;
            rom[2256] = 8'hf7 ;
            rom[2257] = 8'h17 ;
            rom[2258] = 8'hf5 ;
            rom[2259] = 8'hf6 ;
            rom[2260] = 8'h06 ;
            rom[2261] = 8'hfd ;
            rom[2262] = 8'h14 ;
            rom[2263] = 8'hdd ;
            rom[2264] = 8'hfb ;
            rom[2265] = 8'h17 ;
            rom[2266] = 8'h04 ;
            rom[2267] = 8'hd2 ;
            rom[2268] = 8'h01 ;
            rom[2269] = 8'he4 ;
            rom[2270] = 8'hf2 ;
            rom[2271] = 8'hd1 ;
            rom[2272] = 8'h08 ;
            rom[2273] = 8'h0b ;
            rom[2274] = 8'h0a ;
            rom[2275] = 8'h02 ;
            rom[2276] = 8'h01 ;
            rom[2277] = 8'h07 ;
            rom[2278] = 8'h19 ;
            rom[2279] = 8'hf4 ;
            rom[2280] = 8'hdf ;
            rom[2281] = 8'h03 ;
            rom[2282] = 8'hc1 ;
            rom[2283] = 8'h07 ;
            rom[2284] = 8'h21 ;
            rom[2285] = 8'he9 ;
            rom[2286] = 8'h13 ;
            rom[2287] = 8'h0a ;
            rom[2288] = 8'hf7 ;
            rom[2289] = 8'hfa ;
            rom[2290] = 8'h01 ;
            rom[2291] = 8'hfd ;
            rom[2292] = 8'hef ;
            rom[2293] = 8'he4 ;
            rom[2294] = 8'h24 ;
            rom[2295] = 8'hcf ;
            rom[2296] = 8'h01 ;
            rom[2297] = 8'h0b ;
            rom[2298] = 8'hea ;
            rom[2299] = 8'h02 ;
            rom[2300] = 8'hf2 ;
            rom[2301] = 8'hed ;
            rom[2302] = 8'h08 ;
            rom[2303] = 8'hea ;
            rom[2304] = 8'h25 ;
            rom[2305] = 8'hf6 ;
            rom[2306] = 8'he7 ;
            rom[2307] = 8'hf4 ;
            rom[2308] = 8'h01 ;
            rom[2309] = 8'h02 ;
            rom[2310] = 8'h19 ;
            rom[2311] = 8'h16 ;
            rom[2312] = 8'h01 ;
            rom[2313] = 8'h09 ;
            rom[2314] = 8'hef ;
            rom[2315] = 8'hf6 ;
            rom[2316] = 8'he6 ;
            rom[2317] = 8'hf6 ;
            rom[2318] = 8'hf1 ;
            rom[2319] = 8'h0c ;
            rom[2320] = 8'h1e ;
            rom[2321] = 8'h05 ;
            rom[2322] = 8'hec ;
            rom[2323] = 8'hf6 ;
            rom[2324] = 8'h0f ;
            rom[2325] = 8'he4 ;
            rom[2326] = 8'h0a ;
            rom[2327] = 8'h25 ;
            rom[2328] = 8'h07 ;
            rom[2329] = 8'h06 ;
            rom[2330] = 8'h03 ;
            rom[2331] = 8'h0a ;
            rom[2332] = 8'h0a ;
            rom[2333] = 8'hfc ;
            rom[2334] = 8'hdb ;
            rom[2335] = 8'h19 ;
            rom[2336] = 8'h0a ;
            rom[2337] = 8'h1c ;
            rom[2338] = 8'h02 ;
            rom[2339] = 8'hfa ;
            rom[2340] = 8'h13 ;
            rom[2341] = 8'hfb ;
            rom[2342] = 8'hf5 ;
            rom[2343] = 8'hf0 ;
            rom[2344] = 8'h1a ;
            rom[2345] = 8'he1 ;
            rom[2346] = 8'hec ;
            rom[2347] = 8'h01 ;
            rom[2348] = 8'h02 ;
            rom[2349] = 8'h0b ;
            rom[2350] = 8'hee ;
            rom[2351] = 8'hff ;
            rom[2352] = 8'hf1 ;
            rom[2353] = 8'h10 ;
            rom[2354] = 8'h12 ;
            rom[2355] = 8'hf9 ;
            rom[2356] = 8'h10 ;
            rom[2357] = 8'hcb ;
            rom[2358] = 8'hf0 ;
            rom[2359] = 8'hf4 ;
            rom[2360] = 8'h0c ;
            rom[2361] = 8'hfb ;
            rom[2362] = 8'hfc ;
            rom[2363] = 8'h0a ;
            rom[2364] = 8'hfd ;
            rom[2365] = 8'hf5 ;
            rom[2366] = 8'hf0 ;
            rom[2367] = 8'hfe ;
            rom[2368] = 8'hfe ;
            rom[2369] = 8'he9 ;
            rom[2370] = 8'h04 ;
            rom[2371] = 8'h11 ;
            rom[2372] = 8'hf6 ;
            rom[2373] = 8'h02 ;
            rom[2374] = 8'hff ;
            rom[2375] = 8'hf8 ;
            rom[2376] = 8'hf3 ;
            rom[2377] = 8'hd8 ;
            rom[2378] = 8'hf6 ;
            rom[2379] = 8'h01 ;
            rom[2380] = 8'h07 ;
            rom[2381] = 8'hea ;
            rom[2382] = 8'hfd ;
            rom[2383] = 8'h12 ;
            rom[2384] = 8'h00 ;
            rom[2385] = 8'h17 ;
            rom[2386] = 8'hfa ;
            rom[2387] = 8'hf2 ;
            rom[2388] = 8'h07 ;
            rom[2389] = 8'h19 ;
            rom[2390] = 8'h0b ;
            rom[2391] = 8'he0 ;
            rom[2392] = 8'hf7 ;
            rom[2393] = 8'h25 ;
            rom[2394] = 8'h0c ;
            rom[2395] = 8'h11 ;
            rom[2396] = 8'h10 ;
            rom[2397] = 8'h10 ;
            rom[2398] = 8'h12 ;
            rom[2399] = 8'h02 ;
            rom[2400] = 8'h17 ;
            rom[2401] = 8'h12 ;
            rom[2402] = 8'hab ;
            rom[2403] = 8'hfe ;
            rom[2404] = 8'hef ;
            rom[2405] = 8'h1c ;
            rom[2406] = 8'hf9 ;
            rom[2407] = 8'h11 ;
            rom[2408] = 8'hfa ;
            rom[2409] = 8'h06 ;
            rom[2410] = 8'h0f ;
            rom[2411] = 8'ha2 ;
            rom[2412] = 8'hff ;
            rom[2413] = 8'hf3 ;
            rom[2414] = 8'hfc ;
            rom[2415] = 8'hf2 ;
            rom[2416] = 8'h0a ;
            rom[2417] = 8'he8 ;
            rom[2418] = 8'hfc ;
            rom[2419] = 8'hfa ;
            rom[2420] = 8'hfa ;
            rom[2421] = 8'hf0 ;
            rom[2422] = 8'h06 ;
            rom[2423] = 8'h0f ;
            rom[2424] = 8'hf0 ;
            rom[2425] = 8'h02 ;
            rom[2426] = 8'h0c ;
            rom[2427] = 8'h04 ;
            rom[2428] = 8'h15 ;
            rom[2429] = 8'hff ;
            rom[2430] = 8'h08 ;
            rom[2431] = 8'h32 ;
            rom[2432] = 8'h05 ;
            rom[2433] = 8'h08 ;
            rom[2434] = 8'h08 ;
            rom[2435] = 8'h17 ;
            rom[2436] = 8'h07 ;
            rom[2437] = 8'hf7 ;
            rom[2438] = 8'hf7 ;
            rom[2439] = 8'h11 ;
            rom[2440] = 8'h0b ;
            rom[2441] = 8'hfc ;
            rom[2442] = 8'hf9 ;
            rom[2443] = 8'hf9 ;
            rom[2444] = 8'hf0 ;
            rom[2445] = 8'he4 ;
            rom[2446] = 8'h10 ;
            rom[2447] = 8'h15 ;
            rom[2448] = 8'h00 ;
            rom[2449] = 8'hf1 ;
            rom[2450] = 8'h1d ;
            rom[2451] = 8'h10 ;
            rom[2452] = 8'hfe ;
            rom[2453] = 8'h06 ;
            rom[2454] = 8'h19 ;
            rom[2455] = 8'hf5 ;
            rom[2456] = 8'hdb ;
            rom[2457] = 8'h01 ;
            rom[2458] = 8'hf3 ;
            rom[2459] = 8'hff ;
            rom[2460] = 8'hce ;
            rom[2461] = 8'h20 ;
            rom[2462] = 8'he6 ;
            rom[2463] = 8'hd8 ;
            rom[2464] = 8'h09 ;
            rom[2465] = 8'h0f ;
            rom[2466] = 8'h09 ;
            rom[2467] = 8'he5 ;
            rom[2468] = 8'hfa ;
            rom[2469] = 8'h11 ;
            rom[2470] = 8'h17 ;
            rom[2471] = 8'h00 ;
            rom[2472] = 8'h04 ;
            rom[2473] = 8'h11 ;
            rom[2474] = 8'hfc ;
            rom[2475] = 8'hf4 ;
            rom[2476] = 8'h03 ;
            rom[2477] = 8'he4 ;
            rom[2478] = 8'h07 ;
            rom[2479] = 8'h13 ;
            rom[2480] = 8'hf4 ;
            rom[2481] = 8'hf7 ;
            rom[2482] = 8'hda ;
            rom[2483] = 8'h02 ;
            rom[2484] = 8'h16 ;
            rom[2485] = 8'he5 ;
            rom[2486] = 8'hf7 ;
            rom[2487] = 8'h18 ;
            rom[2488] = 8'he9 ;
            rom[2489] = 8'h19 ;
            rom[2490] = 8'hd4 ;
            rom[2491] = 8'h2a ;
            rom[2492] = 8'hea ;
            rom[2493] = 8'he1 ;
            rom[2494] = 8'h0d ;
            rom[2495] = 8'hce ;
            rom[2496] = 8'h03 ;
            rom[2497] = 8'he5 ;
            rom[2498] = 8'h17 ;
            rom[2499] = 8'hd8 ;
            rom[2500] = 8'hf6 ;
            rom[2501] = 8'h23 ;
            rom[2502] = 8'he2 ;
            rom[2503] = 8'hfe ;
            rom[2504] = 8'h14 ;
            rom[2505] = 8'h00 ;
            rom[2506] = 8'h0b ;
            rom[2507] = 8'h0d ;
            rom[2508] = 8'h19 ;
            rom[2509] = 8'h06 ;
            rom[2510] = 8'h0d ;
            rom[2511] = 8'hec ;
            rom[2512] = 8'h0d ;
            rom[2513] = 8'h10 ;
            rom[2514] = 8'hf1 ;
            rom[2515] = 8'hf3 ;
            rom[2516] = 8'h14 ;
            rom[2517] = 8'hcb ;
            rom[2518] = 8'h09 ;
            rom[2519] = 8'hee ;
            rom[2520] = 8'hed ;
            rom[2521] = 8'h14 ;
            rom[2522] = 8'h02 ;
            rom[2523] = 8'hfc ;
            rom[2524] = 8'h16 ;
            rom[2525] = 8'he9 ;
            rom[2526] = 8'hf8 ;
            rom[2527] = 8'h18 ;
            rom[2528] = 8'h22 ;
            rom[2529] = 8'he4 ;
            rom[2530] = 8'h09 ;
            rom[2531] = 8'h16 ;
            rom[2532] = 8'h15 ;
            rom[2533] = 8'h15 ;
            rom[2534] = 8'hff ;
            rom[2535] = 8'h03 ;
            rom[2536] = 8'hf6 ;
            rom[2537] = 8'hfd ;
            rom[2538] = 8'he9 ;
            rom[2539] = 8'hf9 ;
            rom[2540] = 8'h12 ;
            rom[2541] = 8'h0a ;
            rom[2542] = 8'hf9 ;
            rom[2543] = 8'h00 ;
            rom[2544] = 8'hf5 ;
            rom[2545] = 8'h03 ;
            rom[2546] = 8'hff ;
            rom[2547] = 8'h11 ;
            rom[2548] = 8'h0d ;
            rom[2549] = 8'hf2 ;
            rom[2550] = 8'hef ;
            rom[2551] = 8'he1 ;
            rom[2552] = 8'h1f ;
            rom[2553] = 8'hf6 ;
            rom[2554] = 8'hc4 ;
            rom[2555] = 8'h02 ;
            rom[2556] = 8'h02 ;
            rom[2557] = 8'hcf ;
            rom[2558] = 8'h2f ;
            rom[2559] = 8'hea ;
            rom[2560] = 8'h0b ;
            rom[2561] = 8'h1d ;
            rom[2562] = 8'hcf ;
            rom[2563] = 8'hd8 ;
            rom[2564] = 8'hfc ;
            rom[2565] = 8'h17 ;
            rom[2566] = 8'h00 ;
            rom[2567] = 8'hf7 ;
            rom[2568] = 8'h07 ;
            rom[2569] = 8'hf6 ;
            rom[2570] = 8'he4 ;
            rom[2571] = 8'hfb ;
            rom[2572] = 8'h01 ;
            rom[2573] = 8'he4 ;
            rom[2574] = 8'h0e ;
            rom[2575] = 8'h28 ;
            rom[2576] = 8'h0e ;
            rom[2577] = 8'h00 ;
            rom[2578] = 8'h06 ;
            rom[2579] = 8'hcb ;
            rom[2580] = 8'h08 ;
            rom[2581] = 8'hda ;
            rom[2582] = 8'hfc ;
            rom[2583] = 8'h0b ;
            rom[2584] = 8'h0f ;
            rom[2585] = 8'h0d ;
            rom[2586] = 8'h02 ;
            rom[2587] = 8'he9 ;
            rom[2588] = 8'h04 ;
            rom[2589] = 8'h0f ;
            rom[2590] = 8'h07 ;
            rom[2591] = 8'hc8 ;
            rom[2592] = 8'h14 ;
            rom[2593] = 8'hf2 ;
            rom[2594] = 8'he4 ;
            rom[2595] = 8'h21 ;
            rom[2596] = 8'h10 ;
            rom[2597] = 8'hf5 ;
            rom[2598] = 8'he9 ;
            rom[2599] = 8'h03 ;
            rom[2600] = 8'h07 ;
            rom[2601] = 8'hb5 ;
            rom[2602] = 8'hfb ;
            rom[2603] = 8'hc2 ;
            rom[2604] = 8'h02 ;
            rom[2605] = 8'hff ;
            rom[2606] = 8'h0d ;
            rom[2607] = 8'hf6 ;
            rom[2608] = 8'h02 ;
            rom[2609] = 8'he4 ;
            rom[2610] = 8'h09 ;
            rom[2611] = 8'h0a ;
            rom[2612] = 8'hdd ;
            rom[2613] = 8'h04 ;
            rom[2614] = 8'he0 ;
            rom[2615] = 8'hf0 ;
            rom[2616] = 8'hcd ;
            rom[2617] = 8'hf9 ;
            rom[2618] = 8'hf5 ;
            rom[2619] = 8'h04 ;
            rom[2620] = 8'hf7 ;
            rom[2621] = 8'hea ;
            rom[2622] = 8'hf5 ;
            rom[2623] = 8'hdf ;
            rom[2624] = 8'h18 ;
            rom[2625] = 8'h19 ;
            rom[2626] = 8'hfe ;
            rom[2627] = 8'hd2 ;
            rom[2628] = 8'h0f ;
            rom[2629] = 8'h0e ;
            rom[2630] = 8'hfa ;
            rom[2631] = 8'he4 ;
            rom[2632] = 8'h02 ;
            rom[2633] = 8'h12 ;
            rom[2634] = 8'hf7 ;
            rom[2635] = 8'hec ;
            rom[2636] = 8'hf9 ;
            rom[2637] = 8'hd7 ;
            rom[2638] = 8'hed ;
            rom[2639] = 8'h01 ;
            rom[2640] = 8'h13 ;
            rom[2641] = 8'hfa ;
            rom[2642] = 8'h0d ;
            rom[2643] = 8'hf8 ;
            rom[2644] = 8'hf8 ;
            rom[2645] = 8'he5 ;
            rom[2646] = 8'hf1 ;
            rom[2647] = 8'h1d ;
            rom[2648] = 8'h05 ;
            rom[2649] = 8'h04 ;
            rom[2650] = 8'hd7 ;
            rom[2651] = 8'hfc ;
            rom[2652] = 8'h01 ;
            rom[2653] = 8'h1f ;
            rom[2654] = 8'hef ;
            rom[2655] = 8'hd8 ;
            rom[2656] = 8'h0f ;
            rom[2657] = 8'h12 ;
            rom[2658] = 8'hfe ;
            rom[2659] = 8'h00 ;
            rom[2660] = 8'h1c ;
            rom[2661] = 8'h04 ;
            rom[2662] = 8'hdd ;
            rom[2663] = 8'hf9 ;
            rom[2664] = 8'h03 ;
            rom[2665] = 8'hd0 ;
            rom[2666] = 8'h0c ;
            rom[2667] = 8'he9 ;
            rom[2668] = 8'hf4 ;
            rom[2669] = 8'hf9 ;
            rom[2670] = 8'h19 ;
            rom[2671] = 8'h14 ;
            rom[2672] = 8'h13 ;
            rom[2673] = 8'h01 ;
            rom[2674] = 8'h11 ;
            rom[2675] = 8'h05 ;
            rom[2676] = 8'hed ;
            rom[2677] = 8'hf5 ;
            rom[2678] = 8'hf1 ;
            rom[2679] = 8'he2 ;
            rom[2680] = 8'hdb ;
            rom[2681] = 8'hf2 ;
            rom[2682] = 8'he5 ;
            rom[2683] = 8'h02 ;
            rom[2684] = 8'h1a ;
            rom[2685] = 8'hf3 ;
            rom[2686] = 8'hf3 ;
            rom[2687] = 8'hfb ;
            rom[2688] = 8'hf8 ;
            rom[2689] = 8'hdd ;
            rom[2690] = 8'he1 ;
            rom[2691] = 8'h13 ;
            rom[2692] = 8'hee ;
            rom[2693] = 8'h12 ;
            rom[2694] = 8'h1f ;
            rom[2695] = 8'hc9 ;
            rom[2696] = 8'hfc ;
            rom[2697] = 8'hee ;
            rom[2698] = 8'h0d ;
            rom[2699] = 8'hf9 ;
            rom[2700] = 8'hfb ;
            rom[2701] = 8'h09 ;
            rom[2702] = 8'h24 ;
            rom[2703] = 8'h22 ;
            rom[2704] = 8'hf7 ;
            rom[2705] = 8'hfe ;
            rom[2706] = 8'hee ;
            rom[2707] = 8'h0a ;
            rom[2708] = 8'h07 ;
            rom[2709] = 8'h1e ;
            rom[2710] = 8'hfc ;
            rom[2711] = 8'hef ;
            rom[2712] = 8'h1a ;
            rom[2713] = 8'h0a ;
            rom[2714] = 8'hfe ;
            rom[2715] = 8'hd7 ;
            rom[2716] = 8'h03 ;
            rom[2717] = 8'hee ;
            rom[2718] = 8'h38 ;
            rom[2719] = 8'hea ;
            rom[2720] = 8'h09 ;
            rom[2721] = 8'h22 ;
            rom[2722] = 8'h0f ;
            rom[2723] = 8'hf7 ;
            rom[2724] = 8'hea ;
            rom[2725] = 8'h23 ;
            rom[2726] = 8'hfe ;
            rom[2727] = 8'h00 ;
            rom[2728] = 8'he6 ;
            rom[2729] = 8'h00 ;
            rom[2730] = 8'hfe ;
            rom[2731] = 8'h01 ;
            rom[2732] = 8'h2d ;
            rom[2733] = 8'hf6 ;
            rom[2734] = 8'h16 ;
            rom[2735] = 8'h0a ;
            rom[2736] = 8'he4 ;
            rom[2737] = 8'h10 ;
            rom[2738] = 8'h03 ;
            rom[2739] = 8'h27 ;
            rom[2740] = 8'he7 ;
            rom[2741] = 8'hef ;
            rom[2742] = 8'hf9 ;
            rom[2743] = 8'hb0 ;
            rom[2744] = 8'h09 ;
            rom[2745] = 8'h11 ;
            rom[2746] = 8'hef ;
            rom[2747] = 8'h07 ;
            rom[2748] = 8'h35 ;
            rom[2749] = 8'hfc ;
            rom[2750] = 8'hef ;
            rom[2751] = 8'h25 ;
            rom[2752] = 8'h11 ;
            rom[2753] = 8'h22 ;
            rom[2754] = 8'hea ;
            rom[2755] = 8'heb ;
            rom[2756] = 8'h23 ;
            rom[2757] = 8'h1a ;
            rom[2758] = 8'hea ;
            rom[2759] = 8'hf4 ;
            rom[2760] = 8'h23 ;
            rom[2761] = 8'he9 ;
            rom[2762] = 8'hf3 ;
            rom[2763] = 8'h13 ;
            rom[2764] = 8'h1f ;
            rom[2765] = 8'hf2 ;
            rom[2766] = 8'h16 ;
            rom[2767] = 8'h27 ;
            rom[2768] = 8'h1f ;
            rom[2769] = 8'hee ;
            rom[2770] = 8'h07 ;
            rom[2771] = 8'he5 ;
            rom[2772] = 8'h20 ;
            rom[2773] = 8'hf3 ;
            rom[2774] = 8'h09 ;
            rom[2775] = 8'h06 ;
            rom[2776] = 8'h1a ;
            rom[2777] = 8'h05 ;
            rom[2778] = 8'h0a ;
            rom[2779] = 8'he8 ;
            rom[2780] = 8'he7 ;
            rom[2781] = 8'h18 ;
            rom[2782] = 8'h06 ;
            rom[2783] = 8'he7 ;
            rom[2784] = 8'hfc ;
            rom[2785] = 8'h31 ;
            rom[2786] = 8'hf3 ;
            rom[2787] = 8'h07 ;
            rom[2788] = 8'he2 ;
            rom[2789] = 8'heb ;
            rom[2790] = 8'hf3 ;
            rom[2791] = 8'he0 ;
            rom[2792] = 8'he8 ;
            rom[2793] = 8'hef ;
            rom[2794] = 8'h1f ;
            rom[2795] = 8'hd0 ;
            rom[2796] = 8'h1c ;
            rom[2797] = 8'h04 ;
            rom[2798] = 8'he9 ;
            rom[2799] = 8'h02 ;
            rom[2800] = 8'h0c ;
            rom[2801] = 8'he2 ;
            rom[2802] = 8'h03 ;
            rom[2803] = 8'h19 ;
            rom[2804] = 8'h08 ;
            rom[2805] = 8'h0a ;
            rom[2806] = 8'h0e ;
            rom[2807] = 8'hff ;
            rom[2808] = 8'hf2 ;
            rom[2809] = 8'h23 ;
            rom[2810] = 8'hee ;
            rom[2811] = 8'h04 ;
            rom[2812] = 8'hfd ;
            rom[2813] = 8'h0e ;
            rom[2814] = 8'hfa ;
            rom[2815] = 8'hfd ;
            rom[2816] = 8'h1f ;
            rom[2817] = 8'hfe ;
            rom[2818] = 8'h09 ;
            rom[2819] = 8'hf4 ;
            rom[2820] = 8'hfa ;
            rom[2821] = 8'h0a ;
            rom[2822] = 8'he3 ;
            rom[2823] = 8'h0a ;
            rom[2824] = 8'hdf ;
            rom[2825] = 8'h09 ;
            rom[2826] = 8'hec ;
            rom[2827] = 8'hfe ;
            rom[2828] = 8'h07 ;
            rom[2829] = 8'hfb ;
            rom[2830] = 8'hfb ;
            rom[2831] = 8'h0a ;
            rom[2832] = 8'h0d ;
            rom[2833] = 8'hf9 ;
            rom[2834] = 8'h1e ;
            rom[2835] = 8'hfc ;
            rom[2836] = 8'h01 ;
            rom[2837] = 8'h02 ;
            rom[2838] = 8'h20 ;
            rom[2839] = 8'hfb ;
            rom[2840] = 8'hd8 ;
            rom[2841] = 8'h09 ;
            rom[2842] = 8'hf9 ;
            rom[2843] = 8'hf6 ;
            rom[2844] = 8'he4 ;
            rom[2845] = 8'hfc ;
            rom[2846] = 8'hf7 ;
            rom[2847] = 8'h05 ;
            rom[2848] = 8'h09 ;
            rom[2849] = 8'hf2 ;
            rom[2850] = 8'h0e ;
            rom[2851] = 8'hef ;
            rom[2852] = 8'hf7 ;
            rom[2853] = 8'h06 ;
            rom[2854] = 8'h0d ;
            rom[2855] = 8'h15 ;
            rom[2856] = 8'h0d ;
            rom[2857] = 8'h09 ;
            rom[2858] = 8'he2 ;
            rom[2859] = 8'h04 ;
            rom[2860] = 8'hf8 ;
            rom[2861] = 8'hf4 ;
            rom[2862] = 8'h0f ;
            rom[2863] = 8'h12 ;
            rom[2864] = 8'hfd ;
            rom[2865] = 8'h13 ;
            rom[2866] = 8'hf9 ;
            rom[2867] = 8'h00 ;
            rom[2868] = 8'h04 ;
            rom[2869] = 8'hc6 ;
            rom[2870] = 8'h19 ;
            rom[2871] = 8'h0d ;
            rom[2872] = 8'h0d ;
            rom[2873] = 8'h03 ;
            rom[2874] = 8'hcd ;
            rom[2875] = 8'h1b ;
            rom[2876] = 8'he5 ;
            rom[2877] = 8'hd0 ;
            rom[2878] = 8'h17 ;
            rom[2879] = 8'hd7 ;
            rom[2880] = 8'hfa ;
            rom[2881] = 8'h08 ;
            rom[2882] = 8'h01 ;
            rom[2883] = 8'hfd ;
            rom[2884] = 8'hf1 ;
            rom[2885] = 8'h13 ;
            rom[2886] = 8'h0d ;
            rom[2887] = 8'hfb ;
            rom[2888] = 8'hfc ;
            rom[2889] = 8'hf5 ;
            rom[2890] = 8'h07 ;
            rom[2891] = 8'he1 ;
            rom[2892] = 8'hd8 ;
            rom[2893] = 8'hea ;
            rom[2894] = 8'h0c ;
            rom[2895] = 8'h12 ;
            rom[2896] = 8'h10 ;
            rom[2897] = 8'h1b ;
            rom[2898] = 8'h0c ;
            rom[2899] = 8'hc5 ;
            rom[2900] = 8'h11 ;
            rom[2901] = 8'hf7 ;
            rom[2902] = 8'h23 ;
            rom[2903] = 8'h11 ;
            rom[2904] = 8'h02 ;
            rom[2905] = 8'h15 ;
            rom[2906] = 8'h10 ;
            rom[2907] = 8'he0 ;
            rom[2908] = 8'h0f ;
            rom[2909] = 8'hfc ;
            rom[2910] = 8'h0a ;
            rom[2911] = 8'h07 ;
            rom[2912] = 8'hff ;
            rom[2913] = 8'hf7 ;
            rom[2914] = 8'hee ;
            rom[2915] = 8'hff ;
            rom[2916] = 8'hee ;
            rom[2917] = 8'h0e ;
            rom[2918] = 8'h0e ;
            rom[2919] = 8'h0d ;
            rom[2920] = 8'hfa ;
            rom[2921] = 8'hf5 ;
            rom[2922] = 8'hef ;
            rom[2923] = 8'hf8 ;
            rom[2924] = 8'hdc ;
            rom[2925] = 8'hf3 ;
            rom[2926] = 8'hf8 ;
            rom[2927] = 8'he6 ;
            rom[2928] = 8'h02 ;
            rom[2929] = 8'h04 ;
            rom[2930] = 8'h0e ;
            rom[2931] = 8'he4 ;
            rom[2932] = 8'hf7 ;
            rom[2933] = 8'h08 ;
            rom[2934] = 8'hec ;
            rom[2935] = 8'h0d ;
            rom[2936] = 8'hef ;
            rom[2937] = 8'h17 ;
            rom[2938] = 8'he8 ;
            rom[2939] = 8'hf6 ;
            rom[2940] = 8'hf4 ;
            rom[2941] = 8'h03 ;
            rom[2942] = 8'h01 ;
            rom[2943] = 8'hf7 ;
            rom[2944] = 8'h19 ;
            rom[2945] = 8'h0b ;
            rom[2946] = 8'h1c ;
            rom[2947] = 8'hfe ;
            rom[2948] = 8'hf2 ;
            rom[2949] = 8'he8 ;
            rom[2950] = 8'he6 ;
            rom[2951] = 8'hf3 ;
            rom[2952] = 8'h10 ;
            rom[2953] = 8'h16 ;
            rom[2954] = 8'hef ;
            rom[2955] = 8'h19 ;
            rom[2956] = 8'he8 ;
            rom[2957] = 8'hea ;
            rom[2958] = 8'hfb ;
            rom[2959] = 8'h07 ;
            rom[2960] = 8'h0f ;
            rom[2961] = 8'hee ;
            rom[2962] = 8'h0e ;
            rom[2963] = 8'hdb ;
            rom[2964] = 8'hf5 ;
            rom[2965] = 8'h10 ;
            rom[2966] = 8'h13 ;
            rom[2967] = 8'h1b ;
            rom[2968] = 8'hed ;
            rom[2969] = 8'h03 ;
            rom[2970] = 8'hfe ;
            rom[2971] = 8'h04 ;
            rom[2972] = 8'hfd ;
            rom[2973] = 8'h0e ;
            rom[2974] = 8'h0b ;
            rom[2975] = 8'hf8 ;
            rom[2976] = 8'h21 ;
            rom[2977] = 8'hf8 ;
            rom[2978] = 8'h0b ;
            rom[2979] = 8'h0e ;
            rom[2980] = 8'h00 ;
            rom[2981] = 8'hf5 ;
            rom[2982] = 8'h11 ;
            rom[2983] = 8'h04 ;
            rom[2984] = 8'hdc ;
            rom[2985] = 8'h1e ;
            rom[2986] = 8'hf0 ;
            rom[2987] = 8'hf7 ;
            rom[2988] = 8'hfd ;
            rom[2989] = 8'hfe ;
            rom[2990] = 8'hfb ;
            rom[2991] = 8'he9 ;
            rom[2992] = 8'h16 ;
            rom[2993] = 8'hfc ;
            rom[2994] = 8'h10 ;
            rom[2995] = 8'hf9 ;
            rom[2996] = 8'hfe ;
            rom[2997] = 8'hf2 ;
            rom[2998] = 8'hf7 ;
            rom[2999] = 8'h11 ;
            rom[3000] = 8'hee ;
            rom[3001] = 8'h09 ;
            rom[3002] = 8'hf3 ;
            rom[3003] = 8'he3 ;
            rom[3004] = 8'hfe ;
            rom[3005] = 8'h05 ;
            rom[3006] = 8'h09 ;
            rom[3007] = 8'h0f ;
            rom[3008] = 8'hfd ;
            rom[3009] = 8'h0f ;
            rom[3010] = 8'h0e ;
            rom[3011] = 8'h03 ;
            rom[3012] = 8'h07 ;
            rom[3013] = 8'h00 ;
            rom[3014] = 8'hef ;
            rom[3015] = 8'hfd ;
            rom[3016] = 8'h01 ;
            rom[3017] = 8'h17 ;
            rom[3018] = 8'hef ;
            rom[3019] = 8'hfa ;
            rom[3020] = 8'h1c ;
            rom[3021] = 8'hff ;
            rom[3022] = 8'h14 ;
            rom[3023] = 8'hfb ;
            rom[3024] = 8'h11 ;
            rom[3025] = 8'had ;
            rom[3026] = 8'hf7 ;
            rom[3027] = 8'he0 ;
            rom[3028] = 8'hfd ;
            rom[3029] = 8'hed ;
            rom[3030] = 8'hf2 ;
            rom[3031] = 8'h0d ;
            rom[3032] = 8'h05 ;
            rom[3033] = 8'h08 ;
            rom[3034] = 8'hf3 ;
            rom[3035] = 8'h01 ;
            rom[3036] = 8'h05 ;
            rom[3037] = 8'h06 ;
            rom[3038] = 8'h06 ;
            rom[3039] = 8'h02 ;
            rom[3040] = 8'hfd ;
            rom[3041] = 8'h0f ;
            rom[3042] = 8'h1c ;
            rom[3043] = 8'hf7 ;
            rom[3044] = 8'hf6 ;
            rom[3045] = 8'hff ;
            rom[3046] = 8'hf9 ;
            rom[3047] = 8'h00 ;
            rom[3048] = 8'heb ;
            rom[3049] = 8'h05 ;
            rom[3050] = 8'hf1 ;
            rom[3051] = 8'h05 ;
            rom[3052] = 8'hdd ;
            rom[3053] = 8'hed ;
            rom[3054] = 8'h08 ;
            rom[3055] = 8'h16 ;
            rom[3056] = 8'he0 ;
            rom[3057] = 8'hf5 ;
            rom[3058] = 8'h14 ;
            rom[3059] = 8'h02 ;
            rom[3060] = 8'hee ;
            rom[3061] = 8'hc7 ;
            rom[3062] = 8'h21 ;
            rom[3063] = 8'h13 ;
            rom[3064] = 8'hf5 ;
            rom[3065] = 8'h19 ;
            rom[3066] = 8'he2 ;
            rom[3067] = 8'he5 ;
            rom[3068] = 8'hd5 ;
            rom[3069] = 8'hfb ;
            rom[3070] = 8'hfd ;
            rom[3071] = 8'hfc ;
            rom[3072] = 8'h22 ;
            rom[3073] = 8'hee ;
            rom[3074] = 8'h0e ;
            rom[3075] = 8'h03 ;
            rom[3076] = 8'hfa ;
            rom[3077] = 8'hee ;
            rom[3078] = 8'he3 ;
            rom[3079] = 8'hec ;
            rom[3080] = 8'heb ;
            rom[3081] = 8'h09 ;
            rom[3082] = 8'h06 ;
            rom[3083] = 8'he6 ;
            rom[3084] = 8'h13 ;
            rom[3085] = 8'h01 ;
            rom[3086] = 8'h0c ;
            rom[3087] = 8'h1d ;
            rom[3088] = 8'hed ;
            rom[3089] = 8'h02 ;
            rom[3090] = 8'h07 ;
            rom[3091] = 8'hf8 ;
            rom[3092] = 8'h21 ;
            rom[3093] = 8'h0d ;
            rom[3094] = 8'h25 ;
            rom[3095] = 8'h08 ;
            rom[3096] = 8'hdb ;
            rom[3097] = 8'h05 ;
            rom[3098] = 8'hd1 ;
            rom[3099] = 8'h07 ;
            rom[3100] = 8'hdf ;
            rom[3101] = 8'h1e ;
            rom[3102] = 8'hc1 ;
            rom[3103] = 8'he6 ;
            rom[3104] = 8'h14 ;
            rom[3105] = 8'h16 ;
            rom[3106] = 8'h1c ;
            rom[3107] = 8'hd4 ;
            rom[3108] = 8'hf5 ;
            rom[3109] = 8'hf6 ;
            rom[3110] = 8'h1b ;
            rom[3111] = 8'he7 ;
            rom[3112] = 8'h1b ;
            rom[3113] = 8'h00 ;
            rom[3114] = 8'he1 ;
            rom[3115] = 8'hf0 ;
            rom[3116] = 8'hff ;
            rom[3117] = 8'hf8 ;
            rom[3118] = 8'h1c ;
            rom[3119] = 8'h1d ;
            rom[3120] = 8'h04 ;
            rom[3121] = 8'hfc ;
            rom[3122] = 8'hf1 ;
            rom[3123] = 8'h15 ;
            rom[3124] = 8'h1e ;
            rom[3125] = 8'hb7 ;
            rom[3126] = 8'h00 ;
            rom[3127] = 8'h14 ;
            rom[3128] = 8'hd0 ;
            rom[3129] = 8'h03 ;
            rom[3130] = 8'h01 ;
            rom[3131] = 8'hf5 ;
            rom[3132] = 8'he1 ;
            rom[3133] = 8'hdf ;
            rom[3134] = 8'h15 ;
            rom[3135] = 8'hfb ;
            rom[3136] = 8'hfd ;
            rom[3137] = 8'hf6 ;
            rom[3138] = 8'h0e ;
            rom[3139] = 8'he8 ;
            rom[3140] = 8'h04 ;
            rom[3141] = 8'h10 ;
            rom[3142] = 8'h07 ;
            rom[3143] = 8'h0b ;
            rom[3144] = 8'h0b ;
            rom[3145] = 8'hec ;
            rom[3146] = 8'hee ;
            rom[3147] = 8'hfc ;
            rom[3148] = 8'h23 ;
            rom[3149] = 8'h16 ;
            rom[3150] = 8'he8 ;
            rom[3151] = 8'h02 ;
            rom[3152] = 8'hfa ;
            rom[3153] = 8'h0c ;
            rom[3154] = 8'hd7 ;
            rom[3155] = 8'h05 ;
            rom[3156] = 8'h0f ;
            rom[3157] = 8'hfe ;
            rom[3158] = 8'h15 ;
            rom[3159] = 8'hf7 ;
            rom[3160] = 8'hd9 ;
            rom[3161] = 8'h04 ;
            rom[3162] = 8'h09 ;
            rom[3163] = 8'hed ;
            rom[3164] = 8'h06 ;
            rom[3165] = 8'h00 ;
            rom[3166] = 8'hf9 ;
            rom[3167] = 8'h0a ;
            rom[3168] = 8'h03 ;
            rom[3169] = 8'hea ;
            rom[3170] = 8'h08 ;
            rom[3171] = 8'h14 ;
            rom[3172] = 8'h1a ;
            rom[3173] = 8'h21 ;
            rom[3174] = 8'hf8 ;
            rom[3175] = 8'hff ;
            rom[3176] = 8'h1e ;
            rom[3177] = 8'hc9 ;
            rom[3178] = 8'hf8 ;
            rom[3179] = 8'hf3 ;
            rom[3180] = 8'h21 ;
            rom[3181] = 8'h21 ;
            rom[3182] = 8'h00 ;
            rom[3183] = 8'h0f ;
            rom[3184] = 8'h07 ;
            rom[3185] = 8'hf6 ;
            rom[3186] = 8'hdd ;
            rom[3187] = 8'hef ;
            rom[3188] = 8'h03 ;
            rom[3189] = 8'hf6 ;
            rom[3190] = 8'h02 ;
            rom[3191] = 8'he7 ;
            rom[3192] = 8'h1f ;
            rom[3193] = 8'h11 ;
            rom[3194] = 8'hf4 ;
            rom[3195] = 8'h07 ;
            rom[3196] = 8'h15 ;
            rom[3197] = 8'hf2 ;
            rom[3198] = 8'h13 ;
            rom[3199] = 8'hfe ;
            rom[3200] = 8'h08 ;
            rom[3201] = 8'hf7 ;
            rom[3202] = 8'he4 ;
            rom[3203] = 8'hfe ;
            rom[3204] = 8'h07 ;
            rom[3205] = 8'h0c ;
            rom[3206] = 8'h08 ;
            rom[3207] = 8'hed ;
            rom[3208] = 8'hee ;
            rom[3209] = 8'h08 ;
            rom[3210] = 8'hee ;
            rom[3211] = 8'hf4 ;
            rom[3212] = 8'h03 ;
            rom[3213] = 8'hd8 ;
            rom[3214] = 8'hfb ;
            rom[3215] = 8'hfa ;
            rom[3216] = 8'he8 ;
            rom[3217] = 8'h0f ;
            rom[3218] = 8'hf5 ;
            rom[3219] = 8'h04 ;
            rom[3220] = 8'hfd ;
            rom[3221] = 8'he0 ;
            rom[3222] = 8'h1f ;
            rom[3223] = 8'h17 ;
            rom[3224] = 8'he1 ;
            rom[3225] = 8'hfd ;
            rom[3226] = 8'he8 ;
            rom[3227] = 8'hf8 ;
            rom[3228] = 8'hf9 ;
            rom[3229] = 8'h10 ;
            rom[3230] = 8'hf5 ;
            rom[3231] = 8'he8 ;
            rom[3232] = 8'h04 ;
            rom[3233] = 8'hf5 ;
            rom[3234] = 8'hfa ;
            rom[3235] = 8'hff ;
            rom[3236] = 8'hf2 ;
            rom[3237] = 8'h0f ;
            rom[3238] = 8'h08 ;
            rom[3239] = 8'heb ;
            rom[3240] = 8'h03 ;
            rom[3241] = 8'hfb ;
            rom[3242] = 8'h12 ;
            rom[3243] = 8'h13 ;
            rom[3244] = 8'hfc ;
            rom[3245] = 8'hf8 ;
            rom[3246] = 8'h07 ;
            rom[3247] = 8'hfe ;
            rom[3248] = 8'hf9 ;
            rom[3249] = 8'h05 ;
            rom[3250] = 8'h03 ;
            rom[3251] = 8'hed ;
            rom[3252] = 8'h01 ;
            rom[3253] = 8'hef ;
            rom[3254] = 8'h06 ;
            rom[3255] = 8'h13 ;
            rom[3256] = 8'h02 ;
            rom[3257] = 8'hf9 ;
            rom[3258] = 8'h0c ;
            rom[3259] = 8'h0a ;
            rom[3260] = 8'hdc ;
            rom[3261] = 8'h10 ;
            rom[3262] = 8'hfe ;
            rom[3263] = 8'hcd ;
            rom[3264] = 8'hde ;
            rom[3265] = 8'hf7 ;
            rom[3266] = 8'heb ;
            rom[3267] = 8'hf9 ;
            rom[3268] = 8'hfb ;
            rom[3269] = 8'hf8 ;
            rom[3270] = 8'h10 ;
            rom[3271] = 8'h06 ;
            rom[3272] = 8'h22 ;
            rom[3273] = 8'hf0 ;
            rom[3274] = 8'hbd ;
            rom[3275] = 8'hfc ;
            rom[3276] = 8'hfd ;
            rom[3277] = 8'hdd ;
            rom[3278] = 8'hfb ;
            rom[3279] = 8'hfb ;
            rom[3280] = 8'h11 ;
            rom[3281] = 8'h19 ;
            rom[3282] = 8'h12 ;
            rom[3283] = 8'hf4 ;
            rom[3284] = 8'h16 ;
            rom[3285] = 8'h02 ;
            rom[3286] = 8'hf3 ;
            rom[3287] = 8'hfe ;
            rom[3288] = 8'h1b ;
            rom[3289] = 8'h19 ;
            rom[3290] = 8'h04 ;
            rom[3291] = 8'h00 ;
            rom[3292] = 8'hfe ;
            rom[3293] = 8'h02 ;
            rom[3294] = 8'h11 ;
            rom[3295] = 8'hc9 ;
            rom[3296] = 8'h00 ;
            rom[3297] = 8'h0a ;
            rom[3298] = 8'hfe ;
            rom[3299] = 8'hf3 ;
            rom[3300] = 8'hdf ;
            rom[3301] = 8'hf6 ;
            rom[3302] = 8'hd9 ;
            rom[3303] = 8'h09 ;
            rom[3304] = 8'h29 ;
            rom[3305] = 8'hd3 ;
            rom[3306] = 8'hf2 ;
            rom[3307] = 8'h15 ;
            rom[3308] = 8'hee ;
            rom[3309] = 8'hfe ;
            rom[3310] = 8'hec ;
            rom[3311] = 8'h0f ;
            rom[3312] = 8'h03 ;
            rom[3313] = 8'hee ;
            rom[3314] = 8'h1d ;
            rom[3315] = 8'h01 ;
            rom[3316] = 8'h0e ;
            rom[3317] = 8'h09 ;
            rom[3318] = 8'hd3 ;
            rom[3319] = 8'hfb ;
            rom[3320] = 8'he3 ;
            rom[3321] = 8'h0c ;
            rom[3322] = 8'hfc ;
            rom[3323] = 8'h0b ;
            rom[3324] = 8'h0a ;
            rom[3325] = 8'h17 ;
            rom[3326] = 8'hf8 ;
            rom[3327] = 8'h20 ;
            rom[3328] = 8'h29 ;
            rom[3329] = 8'h04 ;
            rom[3330] = 8'h0b ;
            rom[3331] = 8'h07 ;
            rom[3332] = 8'h03 ;
            rom[3333] = 8'h01 ;
            rom[3334] = 8'hf4 ;
            rom[3335] = 8'hf9 ;
            rom[3336] = 8'hf6 ;
            rom[3337] = 8'h1d ;
            rom[3338] = 8'hf0 ;
            rom[3339] = 8'hf4 ;
            rom[3340] = 8'hf6 ;
            rom[3341] = 8'hb6 ;
            rom[3342] = 8'he3 ;
            rom[3343] = 8'h04 ;
            rom[3344] = 8'hf7 ;
            rom[3345] = 8'h21 ;
            rom[3346] = 8'hfb ;
            rom[3347] = 8'h09 ;
            rom[3348] = 8'h10 ;
            rom[3349] = 8'h02 ;
            rom[3350] = 8'h15 ;
            rom[3351] = 8'h06 ;
            rom[3352] = 8'he0 ;
            rom[3353] = 8'h01 ;
            rom[3354] = 8'hde ;
            rom[3355] = 8'h00 ;
            rom[3356] = 8'hf3 ;
            rom[3357] = 8'h10 ;
            rom[3358] = 8'hb9 ;
            rom[3359] = 8'he7 ;
            rom[3360] = 8'h10 ;
            rom[3361] = 8'hfa ;
            rom[3362] = 8'hf5 ;
            rom[3363] = 8'hf4 ;
            rom[3364] = 8'h11 ;
            rom[3365] = 8'hf9 ;
            rom[3366] = 8'h10 ;
            rom[3367] = 8'h07 ;
            rom[3368] = 8'h11 ;
            rom[3369] = 8'hd7 ;
            rom[3370] = 8'h05 ;
            rom[3371] = 8'h01 ;
            rom[3372] = 8'hff ;
            rom[3373] = 8'h08 ;
            rom[3374] = 8'h1c ;
            rom[3375] = 8'h02 ;
            rom[3376] = 8'h25 ;
            rom[3377] = 8'h07 ;
            rom[3378] = 8'h01 ;
            rom[3379] = 8'h0f ;
            rom[3380] = 8'h0d ;
            rom[3381] = 8'he9 ;
            rom[3382] = 8'hea ;
            rom[3383] = 8'hff ;
            rom[3384] = 8'h16 ;
            rom[3385] = 8'hc7 ;
            rom[3386] = 8'h0e ;
            rom[3387] = 8'hfe ;
            rom[3388] = 8'h11 ;
            rom[3389] = 8'h02 ;
            rom[3390] = 8'hde ;
            rom[3391] = 8'he1 ;
            rom[3392] = 8'h0c ;
            rom[3393] = 8'he8 ;
            rom[3394] = 8'hf0 ;
            rom[3395] = 8'hff ;
            rom[3396] = 8'h1c ;
            rom[3397] = 8'hde ;
            rom[3398] = 8'hd7 ;
            rom[3399] = 8'hf8 ;
            rom[3400] = 8'hf9 ;
            rom[3401] = 8'hef ;
            rom[3402] = 8'he8 ;
            rom[3403] = 8'h0e ;
            rom[3404] = 8'h0c ;
            rom[3405] = 8'hf3 ;
            rom[3406] = 8'h21 ;
            rom[3407] = 8'h19 ;
            rom[3408] = 8'h14 ;
            rom[3409] = 8'h14 ;
            rom[3410] = 8'hf4 ;
            rom[3411] = 8'h15 ;
            rom[3412] = 8'h0d ;
            rom[3413] = 8'h02 ;
            rom[3414] = 8'h17 ;
            rom[3415] = 8'h1b ;
            rom[3416] = 8'h08 ;
            rom[3417] = 8'h19 ;
            rom[3418] = 8'hf5 ;
            rom[3419] = 8'h08 ;
            rom[3420] = 8'hf7 ;
            rom[3421] = 8'hf4 ;
            rom[3422] = 8'h02 ;
            rom[3423] = 8'hde ;
            rom[3424] = 8'h19 ;
            rom[3425] = 8'h1d ;
            rom[3426] = 8'hee ;
            rom[3427] = 8'h0d ;
            rom[3428] = 8'hdc ;
            rom[3429] = 8'hf5 ;
            rom[3430] = 8'hf9 ;
            rom[3431] = 8'hf0 ;
            rom[3432] = 8'hf5 ;
            rom[3433] = 8'h0e ;
            rom[3434] = 8'hfe ;
            rom[3435] = 8'hd1 ;
            rom[3436] = 8'hfd ;
            rom[3437] = 8'hef ;
            rom[3438] = 8'hf5 ;
            rom[3439] = 8'h14 ;
            rom[3440] = 8'hfa ;
            rom[3441] = 8'hfa ;
            rom[3442] = 8'h01 ;
            rom[3443] = 8'hdc ;
            rom[3444] = 8'h05 ;
            rom[3445] = 8'hdb ;
            rom[3446] = 8'h03 ;
            rom[3447] = 8'hfb ;
            rom[3448] = 8'hc8 ;
            rom[3449] = 8'he9 ;
            rom[3450] = 8'h10 ;
            rom[3451] = 8'h19 ;
            rom[3452] = 8'hff ;
            rom[3453] = 8'h05 ;
            rom[3454] = 8'hf1 ;
            rom[3455] = 8'h19 ;
            rom[3456] = 8'h07 ;
            rom[3457] = 8'he6 ;
            rom[3458] = 8'h04 ;
            rom[3459] = 8'hec ;
            rom[3460] = 8'hf9 ;
            rom[3461] = 8'h0f ;
            rom[3462] = 8'hf6 ;
            rom[3463] = 8'he0 ;
            rom[3464] = 8'he9 ;
            rom[3465] = 8'hf7 ;
            rom[3466] = 8'hfd ;
            rom[3467] = 8'hff ;
            rom[3468] = 8'hf2 ;
            rom[3469] = 8'hf0 ;
            rom[3470] = 8'he9 ;
            rom[3471] = 8'h0b ;
            rom[3472] = 8'h02 ;
            rom[3473] = 8'h0b ;
            rom[3474] = 8'hf2 ;
            rom[3475] = 8'he7 ;
            rom[3476] = 8'h24 ;
            rom[3477] = 8'he9 ;
            rom[3478] = 8'h16 ;
            rom[3479] = 8'hfe ;
            rom[3480] = 8'he3 ;
            rom[3481] = 8'h12 ;
            rom[3482] = 8'h05 ;
            rom[3483] = 8'h17 ;
            rom[3484] = 8'h11 ;
            rom[3485] = 8'h0d ;
            rom[3486] = 8'h09 ;
            rom[3487] = 8'h03 ;
            rom[3488] = 8'h14 ;
            rom[3489] = 8'h07 ;
            rom[3490] = 8'hc0 ;
            rom[3491] = 8'h03 ;
            rom[3492] = 8'h08 ;
            rom[3493] = 8'h05 ;
            rom[3494] = 8'hdf ;
            rom[3495] = 8'h18 ;
            rom[3496] = 8'h0b ;
            rom[3497] = 8'h06 ;
            rom[3498] = 8'h1a ;
            rom[3499] = 8'hf1 ;
            rom[3500] = 8'hdf ;
            rom[3501] = 8'hf7 ;
            rom[3502] = 8'hfa ;
            rom[3503] = 8'hfd ;
            rom[3504] = 8'hfe ;
            rom[3505] = 8'hd0 ;
            rom[3506] = 8'hf0 ;
            rom[3507] = 8'hf0 ;
            rom[3508] = 8'heb ;
            rom[3509] = 8'h00 ;
            rom[3510] = 8'he6 ;
            rom[3511] = 8'h04 ;
            rom[3512] = 8'h00 ;
            rom[3513] = 8'h0a ;
            rom[3514] = 8'hec ;
            rom[3515] = 8'hfe ;
            rom[3516] = 8'hff ;
            rom[3517] = 8'hf8 ;
            rom[3518] = 8'h05 ;
            rom[3519] = 8'h08 ;
            rom[3520] = 8'heb ;
            rom[3521] = 8'he7 ;
            rom[3522] = 8'he1 ;
            rom[3523] = 8'hea ;
            rom[3524] = 8'hfb ;
            rom[3525] = 8'he9 ;
            rom[3526] = 8'hfa ;
            rom[3527] = 8'h00 ;
            rom[3528] = 8'h12 ;
            rom[3529] = 8'h03 ;
            rom[3530] = 8'hdf ;
            rom[3531] = 8'h11 ;
            rom[3532] = 8'hf0 ;
            rom[3533] = 8'hf8 ;
            rom[3534] = 8'h24 ;
            rom[3535] = 8'h0c ;
            rom[3536] = 8'h21 ;
            rom[3537] = 8'h07 ;
            rom[3538] = 8'hd9 ;
            rom[3539] = 8'h17 ;
            rom[3540] = 8'hfc ;
            rom[3541] = 8'hed ;
            rom[3542] = 8'h0a ;
            rom[3543] = 8'h1f ;
            rom[3544] = 8'h23 ;
            rom[3545] = 8'h0b ;
            rom[3546] = 8'hf5 ;
            rom[3547] = 8'h17 ;
            rom[3548] = 8'hf1 ;
            rom[3549] = 8'hf3 ;
            rom[3550] = 8'h16 ;
            rom[3551] = 8'hf3 ;
            rom[3552] = 8'h12 ;
            rom[3553] = 8'h0c ;
            rom[3554] = 8'hf0 ;
            rom[3555] = 8'hf8 ;
            rom[3556] = 8'hf0 ;
            rom[3557] = 8'hec ;
            rom[3558] = 8'h05 ;
            rom[3559] = 8'hf9 ;
            rom[3560] = 8'hf5 ;
            rom[3561] = 8'h08 ;
            rom[3562] = 8'hff ;
            rom[3563] = 8'hdb ;
            rom[3564] = 8'h11 ;
            rom[3565] = 8'h0f ;
            rom[3566] = 8'he9 ;
            rom[3567] = 8'hf4 ;
            rom[3568] = 8'hef ;
            rom[3569] = 8'h10 ;
            rom[3570] = 8'h03 ;
            rom[3571] = 8'hf0 ;
            rom[3572] = 8'hfd ;
            rom[3573] = 8'hcb ;
            rom[3574] = 8'h0f ;
            rom[3575] = 8'h02 ;
            rom[3576] = 8'hc2 ;
            rom[3577] = 8'hcf ;
            rom[3578] = 8'h12 ;
            rom[3579] = 8'h25 ;
            rom[3580] = 8'hff ;
            rom[3581] = 8'h07 ;
            rom[3582] = 8'h2c ;
            rom[3583] = 8'hef ;
            rom[3584] = 8'h03 ;
            rom[3585] = 8'hcf ;
            rom[3586] = 8'h15 ;
            rom[3587] = 8'hdb ;
            rom[3588] = 8'hf5 ;
            rom[3589] = 8'h0e ;
            rom[3590] = 8'h0e ;
            rom[3591] = 8'h0b ;
            rom[3592] = 8'hec ;
            rom[3593] = 8'hf5 ;
            rom[3594] = 8'he1 ;
            rom[3595] = 8'hf5 ;
            rom[3596] = 8'hfd ;
            rom[3597] = 8'hea ;
            rom[3598] = 8'hd1 ;
            rom[3599] = 8'h11 ;
            rom[3600] = 8'h09 ;
            rom[3601] = 8'h0b ;
            rom[3602] = 8'hed ;
            rom[3603] = 8'h01 ;
            rom[3604] = 8'h1b ;
            rom[3605] = 8'he9 ;
            rom[3606] = 8'h14 ;
            rom[3607] = 8'h01 ;
            rom[3608] = 8'hf4 ;
            rom[3609] = 8'h06 ;
            rom[3610] = 8'hf3 ;
            rom[3611] = 8'h04 ;
            rom[3612] = 8'h21 ;
            rom[3613] = 8'hff ;
            rom[3614] = 8'hed ;
            rom[3615] = 8'hea ;
            rom[3616] = 8'h16 ;
            rom[3617] = 8'he2 ;
            rom[3618] = 8'hf7 ;
            rom[3619] = 8'h15 ;
            rom[3620] = 8'hfe ;
            rom[3621] = 8'h1c ;
            rom[3622] = 8'hf3 ;
            rom[3623] = 8'h07 ;
            rom[3624] = 8'h10 ;
            rom[3625] = 8'hdf ;
            rom[3626] = 8'h05 ;
            rom[3627] = 8'he0 ;
            rom[3628] = 8'hf8 ;
            rom[3629] = 8'hf3 ;
            rom[3630] = 8'h0c ;
            rom[3631] = 8'h11 ;
            rom[3632] = 8'h14 ;
            rom[3633] = 8'h21 ;
            rom[3634] = 8'h18 ;
            rom[3635] = 8'hfe ;
            rom[3636] = 8'h00 ;
            rom[3637] = 8'hd8 ;
            rom[3638] = 8'hec ;
            rom[3639] = 8'hec ;
            rom[3640] = 8'h02 ;
            rom[3641] = 8'hf4 ;
            rom[3642] = 8'hcf ;
            rom[3643] = 8'hfa ;
            rom[3644] = 8'h16 ;
            rom[3645] = 8'he2 ;
            rom[3646] = 8'h08 ;
            rom[3647] = 8'hef ;
            rom[3648] = 8'hea ;
            rom[3649] = 8'hf7 ;
            rom[3650] = 8'hc8 ;
            rom[3651] = 8'hdc ;
            rom[3652] = 8'h07 ;
            rom[3653] = 8'h02 ;
            rom[3654] = 8'h04 ;
            rom[3655] = 8'h06 ;
            rom[3656] = 8'h1c ;
            rom[3657] = 8'hf2 ;
            rom[3658] = 8'h81 ;
            rom[3659] = 8'h04 ;
            rom[3660] = 8'hf1 ;
            rom[3661] = 8'hff ;
            rom[3662] = 8'h00 ;
            rom[3663] = 8'h08 ;
            rom[3664] = 8'h1a ;
            rom[3665] = 8'h0f ;
            rom[3666] = 8'h1f ;
            rom[3667] = 8'hea ;
            rom[3668] = 8'h08 ;
            rom[3669] = 8'h13 ;
            rom[3670] = 8'hfc ;
            rom[3671] = 8'hfe ;
            rom[3672] = 8'hf3 ;
            rom[3673] = 8'h1d ;
            rom[3674] = 8'h1a ;
            rom[3675] = 8'hff ;
            rom[3676] = 8'h12 ;
            rom[3677] = 8'h03 ;
            rom[3678] = 8'h0b ;
            rom[3679] = 8'he4 ;
            rom[3680] = 8'h14 ;
            rom[3681] = 8'h0e ;
            rom[3682] = 8'h08 ;
            rom[3683] = 8'h00 ;
            rom[3684] = 8'he1 ;
            rom[3685] = 8'h09 ;
            rom[3686] = 8'he9 ;
            rom[3687] = 8'h0b ;
            rom[3688] = 8'h0c ;
            rom[3689] = 8'hd9 ;
            rom[3690] = 8'h00 ;
            rom[3691] = 8'hd7 ;
            rom[3692] = 8'hf7 ;
            rom[3693] = 8'h09 ;
            rom[3694] = 8'h03 ;
            rom[3695] = 8'hfb ;
            rom[3696] = 8'h15 ;
            rom[3697] = 8'h0a ;
            rom[3698] = 8'h12 ;
            rom[3699] = 8'h03 ;
            rom[3700] = 8'hf3 ;
            rom[3701] = 8'h11 ;
            rom[3702] = 8'hcd ;
            rom[3703] = 8'hfe ;
            rom[3704] = 8'hda ;
            rom[3705] = 8'h0a ;
            rom[3706] = 8'hfb ;
            rom[3707] = 8'hfe ;
            rom[3708] = 8'h04 ;
            rom[3709] = 8'h17 ;
            rom[3710] = 8'hf1 ;
            rom[3711] = 8'h06 ;
            rom[3712] = 8'hf5 ;
            rom[3713] = 8'h0f ;
            rom[3714] = 8'he1 ;
            rom[3715] = 8'hcc ;
            rom[3716] = 8'h0b ;
            rom[3717] = 8'hee ;
            rom[3718] = 8'h05 ;
            rom[3719] = 8'h02 ;
            rom[3720] = 8'hff ;
            rom[3721] = 8'he7 ;
            rom[3722] = 8'hd4 ;
            rom[3723] = 8'h0d ;
            rom[3724] = 8'h0e ;
            rom[3725] = 8'hf8 ;
            rom[3726] = 8'h0c ;
            rom[3727] = 8'h1d ;
            rom[3728] = 8'h1e ;
            rom[3729] = 8'h06 ;
            rom[3730] = 8'h11 ;
            rom[3731] = 8'hd6 ;
            rom[3732] = 8'h04 ;
            rom[3733] = 8'hde ;
            rom[3734] = 8'h02 ;
            rom[3735] = 8'h13 ;
            rom[3736] = 8'h14 ;
            rom[3737] = 8'h27 ;
            rom[3738] = 8'h04 ;
            rom[3739] = 8'hfc ;
            rom[3740] = 8'h09 ;
            rom[3741] = 8'h07 ;
            rom[3742] = 8'hf5 ;
            rom[3743] = 8'hed ;
            rom[3744] = 8'h10 ;
            rom[3745] = 8'hfe ;
            rom[3746] = 8'hd5 ;
            rom[3747] = 8'hfc ;
            rom[3748] = 8'he2 ;
            rom[3749] = 8'hf3 ;
            rom[3750] = 8'he9 ;
            rom[3751] = 8'h05 ;
            rom[3752] = 8'h0b ;
            rom[3753] = 8'hea ;
            rom[3754] = 8'h15 ;
            rom[3755] = 8'h98 ;
            rom[3756] = 8'hf6 ;
            rom[3757] = 8'h0f ;
            rom[3758] = 8'h0d ;
            rom[3759] = 8'hff ;
            rom[3760] = 8'h04 ;
            rom[3761] = 8'hd0 ;
            rom[3762] = 8'h09 ;
            rom[3763] = 8'hf8 ;
            rom[3764] = 8'hdc ;
            rom[3765] = 8'h0f ;
            rom[3766] = 8'hf0 ;
            rom[3767] = 8'h16 ;
            rom[3768] = 8'hda ;
            rom[3769] = 8'h1c ;
            rom[3770] = 8'hf7 ;
            rom[3771] = 8'h1b ;
            rom[3772] = 8'hff ;
            rom[3773] = 8'hf7 ;
            rom[3774] = 8'h0e ;
            rom[3775] = 8'h0a ;
            rom[3776] = 8'hed ;
            rom[3777] = 8'hec ;
            rom[3778] = 8'h00 ;
            rom[3779] = 8'he1 ;
            rom[3780] = 8'h05 ;
            rom[3781] = 8'hcc ;
            rom[3782] = 8'hf4 ;
            rom[3783] = 8'hf9 ;
            rom[3784] = 8'hff ;
            rom[3785] = 8'hf2 ;
            rom[3786] = 8'hc4 ;
            rom[3787] = 8'h09 ;
            rom[3788] = 8'hf5 ;
            rom[3789] = 8'h02 ;
            rom[3790] = 8'h08 ;
            rom[3791] = 8'h1b ;
            rom[3792] = 8'h13 ;
            rom[3793] = 8'h1f ;
            rom[3794] = 8'hf9 ;
            rom[3795] = 8'h0c ;
            rom[3796] = 8'h22 ;
            rom[3797] = 8'h0a ;
            rom[3798] = 8'h0e ;
            rom[3799] = 8'h0c ;
            rom[3800] = 8'h03 ;
            rom[3801] = 8'h05 ;
            rom[3802] = 8'h1b ;
            rom[3803] = 8'h09 ;
            rom[3804] = 8'h17 ;
            rom[3805] = 8'hf5 ;
            rom[3806] = 8'h08 ;
            rom[3807] = 8'he0 ;
            rom[3808] = 8'h17 ;
            rom[3809] = 8'h09 ;
            rom[3810] = 8'hd8 ;
            rom[3811] = 8'h03 ;
            rom[3812] = 8'hef ;
            rom[3813] = 8'h18 ;
            rom[3814] = 8'hfd ;
            rom[3815] = 8'hfb ;
            rom[3816] = 8'h04 ;
            rom[3817] = 8'hf7 ;
            rom[3818] = 8'h15 ;
            rom[3819] = 8'hd5 ;
            rom[3820] = 8'hf8 ;
            rom[3821] = 8'h15 ;
            rom[3822] = 8'hfe ;
            rom[3823] = 8'h00 ;
            rom[3824] = 8'hff ;
            rom[3825] = 8'heb ;
            rom[3826] = 8'h0f ;
            rom[3827] = 8'he8 ;
            rom[3828] = 8'h0a ;
            rom[3829] = 8'he4 ;
            rom[3830] = 8'h13 ;
            rom[3831] = 8'hee ;
            rom[3832] = 8'hd2 ;
            rom[3833] = 8'h07 ;
            rom[3834] = 8'h07 ;
            rom[3835] = 8'h06 ;
            rom[3836] = 8'h0d ;
            rom[3837] = 8'h15 ;
            rom[3838] = 8'h0e ;
            rom[3839] = 8'h02 ;
            rom[3840] = 8'h0b ;
            rom[3841] = 8'hfb ;
            rom[3842] = 8'h04 ;
            rom[3843] = 8'h1e ;
            rom[3844] = 8'h07 ;
            rom[3845] = 8'hee ;
            rom[3846] = 8'hf0 ;
            rom[3847] = 8'h03 ;
            rom[3848] = 8'h0b ;
            rom[3849] = 8'h03 ;
            rom[3850] = 8'hea ;
            rom[3851] = 8'h09 ;
            rom[3852] = 8'hd3 ;
            rom[3853] = 8'hd3 ;
            rom[3854] = 8'h01 ;
            rom[3855] = 8'h00 ;
            rom[3856] = 8'hf9 ;
            rom[3857] = 8'h25 ;
            rom[3858] = 8'hf1 ;
            rom[3859] = 8'hfa ;
            rom[3860] = 8'h07 ;
            rom[3861] = 8'h0b ;
            rom[3862] = 8'h22 ;
            rom[3863] = 8'h04 ;
            rom[3864] = 8'hfd ;
            rom[3865] = 8'h2e ;
            rom[3866] = 8'hef ;
            rom[3867] = 8'h0d ;
            rom[3868] = 8'hf3 ;
            rom[3869] = 8'h0c ;
            rom[3870] = 8'hea ;
            rom[3871] = 8'hee ;
            rom[3872] = 8'h1c ;
            rom[3873] = 8'h0c ;
            rom[3874] = 8'h03 ;
            rom[3875] = 8'h0a ;
            rom[3876] = 8'he6 ;
            rom[3877] = 8'hd2 ;
            rom[3878] = 8'h0f ;
            rom[3879] = 8'he9 ;
            rom[3880] = 8'hd1 ;
            rom[3881] = 8'h08 ;
            rom[3882] = 8'hfd ;
            rom[3883] = 8'h04 ;
            rom[3884] = 8'he7 ;
            rom[3885] = 8'h16 ;
            rom[3886] = 8'h25 ;
            rom[3887] = 8'hee ;
            rom[3888] = 8'h16 ;
            rom[3889] = 8'hf1 ;
            rom[3890] = 8'h10 ;
            rom[3891] = 8'hdd ;
            rom[3892] = 8'h07 ;
            rom[3893] = 8'hd5 ;
            rom[3894] = 8'heb ;
            rom[3895] = 8'h0a ;
            rom[3896] = 8'hd8 ;
            rom[3897] = 8'hde ;
            rom[3898] = 8'h0a ;
            rom[3899] = 8'h03 ;
            rom[3900] = 8'hf8 ;
            rom[3901] = 8'h02 ;
            rom[3902] = 8'hff ;
            rom[3903] = 8'h0c ;
            rom[3904] = 8'h1b ;
            rom[3905] = 8'h19 ;
            rom[3906] = 8'hef ;
            rom[3907] = 8'he9 ;
            rom[3908] = 8'hf6 ;
            rom[3909] = 8'h12 ;
            rom[3910] = 8'hfc ;
            rom[3911] = 8'hdd ;
            rom[3912] = 8'h10 ;
            rom[3913] = 8'hf5 ;
            rom[3914] = 8'h06 ;
            rom[3915] = 8'h08 ;
            rom[3916] = 8'hf5 ;
            rom[3917] = 8'hdf ;
            rom[3918] = 8'h20 ;
            rom[3919] = 8'hf4 ;
            rom[3920] = 8'h0f ;
            rom[3921] = 8'hfb ;
            rom[3922] = 8'hfa ;
            rom[3923] = 8'h0b ;
            rom[3924] = 8'h07 ;
            rom[3925] = 8'he0 ;
            rom[3926] = 8'h08 ;
            rom[3927] = 8'hf3 ;
            rom[3928] = 8'h0e ;
            rom[3929] = 8'hfd ;
            rom[3930] = 8'h11 ;
            rom[3931] = 8'hfa ;
            rom[3932] = 8'h05 ;
            rom[3933] = 8'he5 ;
            rom[3934] = 8'h08 ;
            rom[3935] = 8'hf1 ;
            rom[3936] = 8'h07 ;
            rom[3937] = 8'hf2 ;
            rom[3938] = 8'hfd ;
            rom[3939] = 8'h2f ;
            rom[3940] = 8'h02 ;
            rom[3941] = 8'h00 ;
            rom[3942] = 8'he5 ;
            rom[3943] = 8'hfc ;
            rom[3944] = 8'hf3 ;
            rom[3945] = 8'hd3 ;
            rom[3946] = 8'h14 ;
            rom[3947] = 8'hfe ;
            rom[3948] = 8'hd3 ;
            rom[3949] = 8'h0f ;
            rom[3950] = 8'h02 ;
            rom[3951] = 8'hfa ;
            rom[3952] = 8'h05 ;
            rom[3953] = 8'hfe ;
            rom[3954] = 8'h09 ;
            rom[3955] = 8'h18 ;
            rom[3956] = 8'hc6 ;
            rom[3957] = 8'hfc ;
            rom[3958] = 8'h14 ;
            rom[3959] = 8'h05 ;
            rom[3960] = 8'hf3 ;
            rom[3961] = 8'h02 ;
            rom[3962] = 8'hd5 ;
            rom[3963] = 8'h0b ;
            rom[3964] = 8'h16 ;
            rom[3965] = 8'hfa ;
            rom[3966] = 8'he3 ;
            rom[3967] = 8'hd5 ;
            rom[3968] = 8'he9 ;
            rom[3969] = 8'he6 ;
            rom[3970] = 8'h1a ;
            rom[3971] = 8'heb ;
            rom[3972] = 8'h08 ;
            rom[3973] = 8'h24 ;
            rom[3974] = 8'hc6 ;
            rom[3975] = 8'hdc ;
            rom[3976] = 8'hdc ;
            rom[3977] = 8'h13 ;
            rom[3978] = 8'h07 ;
            rom[3979] = 8'hf4 ;
            rom[3980] = 8'h13 ;
            rom[3981] = 8'hf4 ;
            rom[3982] = 8'hee ;
            rom[3983] = 8'h09 ;
            rom[3984] = 8'hf2 ;
            rom[3985] = 8'h09 ;
            rom[3986] = 8'h14 ;
            rom[3987] = 8'hfc ;
            rom[3988] = 8'h1e ;
            rom[3989] = 8'hca ;
            rom[3990] = 8'h15 ;
            rom[3991] = 8'h17 ;
            rom[3992] = 8'hc8 ;
            rom[3993] = 8'hfc ;
            rom[3994] = 8'he7 ;
            rom[3995] = 8'h01 ;
            rom[3996] = 8'hfc ;
            rom[3997] = 8'h0a ;
            rom[3998] = 8'h0e ;
            rom[3999] = 8'h09 ;
            rom[4000] = 8'h0b ;
            rom[4001] = 8'hfc ;
            rom[4002] = 8'h18 ;
            rom[4003] = 8'hd9 ;
            rom[4004] = 8'h1d ;
            rom[4005] = 8'h18 ;
            rom[4006] = 8'h0b ;
            rom[4007] = 8'h0a ;
            rom[4008] = 8'h13 ;
            rom[4009] = 8'hff ;
            rom[4010] = 8'h05 ;
            rom[4011] = 8'h06 ;
            rom[4012] = 8'hf2 ;
            rom[4013] = 8'hf9 ;
            rom[4014] = 8'he2 ;
            rom[4015] = 8'h00 ;
            rom[4016] = 8'h23 ;
            rom[4017] = 8'he8 ;
            rom[4018] = 8'hf9 ;
            rom[4019] = 8'he2 ;
            rom[4020] = 8'hfe ;
            rom[4021] = 8'hd7 ;
            rom[4022] = 8'h0a ;
            rom[4023] = 8'h18 ;
            rom[4024] = 8'h0c ;
            rom[4025] = 8'h20 ;
            rom[4026] = 8'hcf ;
            rom[4027] = 8'hfd ;
            rom[4028] = 8'hf8 ;
            rom[4029] = 8'hec ;
            rom[4030] = 8'h1c ;
            rom[4031] = 8'hf1 ;
            rom[4032] = 8'h05 ;
            rom[4033] = 8'hfe ;
            rom[4034] = 8'heb ;
            rom[4035] = 8'h00 ;
            rom[4036] = 8'h0c ;
            rom[4037] = 8'h00 ;
            rom[4038] = 8'hf9 ;
            rom[4039] = 8'hfa ;
            rom[4040] = 8'h09 ;
            rom[4041] = 8'hf6 ;
            rom[4042] = 8'h1b ;
            rom[4043] = 8'h0d ;
            rom[4044] = 8'h01 ;
            rom[4045] = 8'h10 ;
            rom[4046] = 8'h14 ;
            rom[4047] = 8'h04 ;
            rom[4048] = 8'h28 ;
            rom[4049] = 8'he3 ;
            rom[4050] = 8'hdd ;
            rom[4051] = 8'hfe ;
            rom[4052] = 8'hf1 ;
            rom[4053] = 8'hd9 ;
            rom[4054] = 8'hee ;
            rom[4055] = 8'hfa ;
            rom[4056] = 8'h1b ;
            rom[4057] = 8'hf8 ;
            rom[4058] = 8'h0a ;
            rom[4059] = 8'h0f ;
            rom[4060] = 8'h05 ;
            rom[4061] = 8'h05 ;
            rom[4062] = 8'hf9 ;
            rom[4063] = 8'he5 ;
            rom[4064] = 8'h04 ;
            rom[4065] = 8'he7 ;
            rom[4066] = 8'h05 ;
            rom[4067] = 8'h19 ;
            rom[4068] = 8'h03 ;
            rom[4069] = 8'heb ;
            rom[4070] = 8'hf4 ;
            rom[4071] = 8'hcd ;
            rom[4072] = 8'hde ;
            rom[4073] = 8'he4 ;
            rom[4074] = 8'h1d ;
            rom[4075] = 8'he2 ;
            rom[4076] = 8'hfe ;
            rom[4077] = 8'hfd ;
            rom[4078] = 8'he0 ;
            rom[4079] = 8'h02 ;
            rom[4080] = 8'he5 ;
            rom[4081] = 8'hd5 ;
            rom[4082] = 8'hf5 ;
            rom[4083] = 8'h18 ;
            rom[4084] = 8'hdd ;
            rom[4085] = 8'h0d ;
            rom[4086] = 8'hfc ;
            rom[4087] = 8'h06 ;
            rom[4088] = 8'hca ;
            rom[4089] = 8'h20 ;
            rom[4090] = 8'hdc ;
            rom[4091] = 8'hfe ;
            rom[4092] = 8'hff ;
            rom[4093] = 8'hf9 ;
            rom[4094] = 8'h19 ;
            rom[4095] = 8'h0f ;
            rom[4096] = 8'h07 ;
            rom[4097] = 8'h0c ;
            rom[4098] = 8'he5 ;
            rom[4099] = 8'h25 ;
            rom[4100] = 8'he5 ;
            rom[4101] = 8'h0d ;
            rom[4102] = 8'hed ;
            rom[4103] = 8'hc3 ;
            rom[4104] = 8'h17 ;
            rom[4105] = 8'hf4 ;
            rom[4106] = 8'h0f ;
            rom[4107] = 8'hf4 ;
            rom[4108] = 8'hcf ;
            rom[4109] = 8'hdd ;
            rom[4110] = 8'h22 ;
            rom[4111] = 8'h09 ;
            rom[4112] = 8'hf4 ;
            rom[4113] = 8'hfa ;
            rom[4114] = 8'hf5 ;
            rom[4115] = 8'he2 ;
            rom[4116] = 8'hf8 ;
            rom[4117] = 8'hdf ;
            rom[4118] = 8'h06 ;
            rom[4119] = 8'h09 ;
            rom[4120] = 8'hf5 ;
            rom[4121] = 8'h0b ;
            rom[4122] = 8'h1d ;
            rom[4123] = 8'h0b ;
            rom[4124] = 8'hdf ;
            rom[4125] = 8'hef ;
            rom[4126] = 8'hef ;
            rom[4127] = 8'he8 ;
            rom[4128] = 8'h07 ;
            rom[4129] = 8'hf1 ;
            rom[4130] = 8'hf0 ;
            rom[4131] = 8'h01 ;
            rom[4132] = 8'h03 ;
            rom[4133] = 8'hff ;
            rom[4134] = 8'h15 ;
            rom[4135] = 8'hf3 ;
            rom[4136] = 8'hee ;
            rom[4137] = 8'he8 ;
            rom[4138] = 8'he1 ;
            rom[4139] = 8'h0d ;
            rom[4140] = 8'hfe ;
            rom[4141] = 8'hea ;
            rom[4142] = 8'h0e ;
            rom[4143] = 8'he6 ;
            rom[4144] = 8'hff ;
            rom[4145] = 8'hfe ;
            rom[4146] = 8'h06 ;
            rom[4147] = 8'h00 ;
            rom[4148] = 8'he9 ;
            rom[4149] = 8'hf0 ;
            rom[4150] = 8'he6 ;
            rom[4151] = 8'hc0 ;
            rom[4152] = 8'h05 ;
            rom[4153] = 8'h01 ;
            rom[4154] = 8'he4 ;
            rom[4155] = 8'he0 ;
            rom[4156] = 8'hff ;
            rom[4157] = 8'hfe ;
            rom[4158] = 8'h01 ;
            rom[4159] = 8'hc9 ;
            rom[4160] = 8'h03 ;
            rom[4161] = 8'hd6 ;
            rom[4162] = 8'hc5 ;
            rom[4163] = 8'hdd ;
            rom[4164] = 8'h17 ;
            rom[4165] = 8'h13 ;
            rom[4166] = 8'hf5 ;
            rom[4167] = 8'hef ;
            rom[4168] = 8'h12 ;
            rom[4169] = 8'h0a ;
            rom[4170] = 8'hef ;
            rom[4171] = 8'hdb ;
            rom[4172] = 8'h15 ;
            rom[4173] = 8'he3 ;
            rom[4174] = 8'hed ;
            rom[4175] = 8'hfa ;
            rom[4176] = 8'h15 ;
            rom[4177] = 8'hfd ;
            rom[4178] = 8'h13 ;
            rom[4179] = 8'hf6 ;
            rom[4180] = 8'hd9 ;
            rom[4181] = 8'hf3 ;
            rom[4182] = 8'h12 ;
            rom[4183] = 8'hf7 ;
            rom[4184] = 8'hf8 ;
            rom[4185] = 8'h0b ;
            rom[4186] = 8'h0f ;
            rom[4187] = 8'hf8 ;
            rom[4188] = 8'hf5 ;
            rom[4189] = 8'h03 ;
            rom[4190] = 8'h17 ;
            rom[4191] = 8'hfc ;
            rom[4192] = 8'h08 ;
            rom[4193] = 8'h0b ;
            rom[4194] = 8'h0c ;
            rom[4195] = 8'he9 ;
            rom[4196] = 8'h1b ;
            rom[4197] = 8'h13 ;
            rom[4198] = 8'h14 ;
            rom[4199] = 8'he6 ;
            rom[4200] = 8'h1c ;
            rom[4201] = 8'he5 ;
            rom[4202] = 8'hf7 ;
            rom[4203] = 8'h13 ;
            rom[4204] = 8'h09 ;
            rom[4205] = 8'he5 ;
            rom[4206] = 8'h14 ;
            rom[4207] = 8'hfa ;
            rom[4208] = 8'h00 ;
            rom[4209] = 8'hea ;
            rom[4210] = 8'h04 ;
            rom[4211] = 8'h13 ;
            rom[4212] = 8'hea ;
            rom[4213] = 8'he0 ;
            rom[4214] = 8'hea ;
            rom[4215] = 8'hfb ;
            rom[4216] = 8'h11 ;
            rom[4217] = 8'h08 ;
            rom[4218] = 8'h08 ;
            rom[4219] = 8'hfe ;
            rom[4220] = 8'h21 ;
            rom[4221] = 8'hfa ;
            rom[4222] = 8'h00 ;
            rom[4223] = 8'he8 ;
            rom[4224] = 8'h03 ;
            rom[4225] = 8'hec ;
            rom[4226] = 8'h19 ;
            rom[4227] = 8'h07 ;
            rom[4228] = 8'hf1 ;
            rom[4229] = 8'hcb ;
            rom[4230] = 8'hdc ;
            rom[4231] = 8'h16 ;
            rom[4232] = 8'hfb ;
            rom[4233] = 8'h1a ;
            rom[4234] = 8'hf8 ;
            rom[4235] = 8'hfe ;
            rom[4236] = 8'h16 ;
            rom[4237] = 8'hfa ;
            rom[4238] = 8'h02 ;
            rom[4239] = 8'h05 ;
            rom[4240] = 8'h09 ;
            rom[4241] = 8'hf6 ;
            rom[4242] = 8'hc0 ;
            rom[4243] = 8'h20 ;
            rom[4244] = 8'hef ;
            rom[4245] = 8'hd1 ;
            rom[4246] = 8'h24 ;
            rom[4247] = 8'hff ;
            rom[4248] = 8'h0b ;
            rom[4249] = 8'hea ;
            rom[4250] = 8'hff ;
            rom[4251] = 8'heb ;
            rom[4252] = 8'h04 ;
            rom[4253] = 8'hf3 ;
            rom[4254] = 8'hdc ;
            rom[4255] = 8'h10 ;
            rom[4256] = 8'hfd ;
            rom[4257] = 8'h0d ;
            rom[4258] = 8'h1a ;
            rom[4259] = 8'h00 ;
            rom[4260] = 8'hee ;
            rom[4261] = 8'heb ;
            rom[4262] = 8'hf7 ;
            rom[4263] = 8'hfd ;
            rom[4264] = 8'hfc ;
            rom[4265] = 8'h0f ;
            rom[4266] = 8'h06 ;
            rom[4267] = 8'hf8 ;
            rom[4268] = 8'hff ;
            rom[4269] = 8'h0d ;
            rom[4270] = 8'h11 ;
            rom[4271] = 8'h0d ;
            rom[4272] = 8'heb ;
            rom[4273] = 8'h08 ;
            rom[4274] = 8'h04 ;
            rom[4275] = 8'h0b ;
            rom[4276] = 8'hfd ;
            rom[4277] = 8'he5 ;
            rom[4278] = 8'hfa ;
            rom[4279] = 8'h14 ;
            rom[4280] = 8'h03 ;
            rom[4281] = 8'h08 ;
            rom[4282] = 8'he5 ;
            rom[4283] = 8'hfa ;
            rom[4284] = 8'h0e ;
            rom[4285] = 8'h02 ;
            rom[4286] = 8'hd9 ;
            rom[4287] = 8'hfe ;
            rom[4288] = 8'h2e ;
            rom[4289] = 8'hef ;
            rom[4290] = 8'h09 ;
            rom[4291] = 8'h03 ;
            rom[4292] = 8'hf9 ;
            rom[4293] = 8'hf8 ;
            rom[4294] = 8'hde ;
            rom[4295] = 8'heb ;
            rom[4296] = 8'hf2 ;
            rom[4297] = 8'hf0 ;
            rom[4298] = 8'h0b ;
            rom[4299] = 8'h13 ;
            rom[4300] = 8'h1c ;
            rom[4301] = 8'he9 ;
            rom[4302] = 8'hfd ;
            rom[4303] = 8'he8 ;
            rom[4304] = 8'hea ;
            rom[4305] = 8'h12 ;
            rom[4306] = 8'h0d ;
            rom[4307] = 8'h06 ;
            rom[4308] = 8'hef ;
            rom[4309] = 8'hfe ;
            rom[4310] = 8'h06 ;
            rom[4311] = 8'hf1 ;
            rom[4312] = 8'h1d ;
            rom[4313] = 8'h0d ;
            rom[4314] = 8'hfa ;
            rom[4315] = 8'hed ;
            rom[4316] = 8'hf8 ;
            rom[4317] = 8'hfb ;
            rom[4318] = 8'hea ;
            rom[4319] = 8'hec ;
            rom[4320] = 8'h14 ;
            rom[4321] = 8'h1a ;
            rom[4322] = 8'h0a ;
            rom[4323] = 8'h11 ;
            rom[4324] = 8'h17 ;
            rom[4325] = 8'h15 ;
            rom[4326] = 8'h12 ;
            rom[4327] = 8'hfd ;
            rom[4328] = 8'hd4 ;
            rom[4329] = 8'h05 ;
            rom[4330] = 8'hea ;
            rom[4331] = 8'h08 ;
            rom[4332] = 8'h17 ;
            rom[4333] = 8'h09 ;
            rom[4334] = 8'h24 ;
            rom[4335] = 8'h18 ;
            rom[4336] = 8'hfe ;
            rom[4337] = 8'hfa ;
            rom[4338] = 8'hff ;
            rom[4339] = 8'h0c ;
            rom[4340] = 8'he1 ;
            rom[4341] = 8'h09 ;
            rom[4342] = 8'h14 ;
            rom[4343] = 8'hcc ;
            rom[4344] = 8'h20 ;
            rom[4345] = 8'hf5 ;
            rom[4346] = 8'hd8 ;
            rom[4347] = 8'h00 ;
            rom[4348] = 8'hfe ;
            rom[4349] = 8'h00 ;
            rom[4350] = 8'hea ;
            rom[4351] = 8'h05 ;
            rom[4352] = 8'h0a ;
            rom[4353] = 8'h0c ;
            rom[4354] = 8'hc8 ;
            rom[4355] = 8'h0c ;
            rom[4356] = 8'h08 ;
            rom[4357] = 8'hed ;
            rom[4358] = 8'h18 ;
            rom[4359] = 8'h1c ;
            rom[4360] = 8'h05 ;
            rom[4361] = 8'h15 ;
            rom[4362] = 8'hdc ;
            rom[4363] = 8'hfe ;
            rom[4364] = 8'hea ;
            rom[4365] = 8'h04 ;
            rom[4366] = 8'hfb ;
            rom[4367] = 8'hfc ;
            rom[4368] = 8'h01 ;
            rom[4369] = 8'h07 ;
            rom[4370] = 8'he6 ;
            rom[4371] = 8'h07 ;
            rom[4372] = 8'h09 ;
            rom[4373] = 8'hd3 ;
            rom[4374] = 8'hfc ;
            rom[4375] = 8'h1b ;
            rom[4376] = 8'hfe ;
            rom[4377] = 8'h06 ;
            rom[4378] = 8'hff ;
            rom[4379] = 8'h1e ;
            rom[4380] = 8'h04 ;
            rom[4381] = 8'h05 ;
            rom[4382] = 8'hed ;
            rom[4383] = 8'hf1 ;
            rom[4384] = 8'hf2 ;
            rom[4385] = 8'h00 ;
            rom[4386] = 8'h01 ;
            rom[4387] = 8'hf9 ;
            rom[4388] = 8'h0d ;
            rom[4389] = 8'hf5 ;
            rom[4390] = 8'hfd ;
            rom[4391] = 8'hed ;
            rom[4392] = 8'h15 ;
            rom[4393] = 8'hfb ;
            rom[4394] = 8'heb ;
            rom[4395] = 8'hfb ;
            rom[4396] = 8'h03 ;
            rom[4397] = 8'hf2 ;
            rom[4398] = 8'h02 ;
            rom[4399] = 8'h0c ;
            rom[4400] = 8'he4 ;
            rom[4401] = 8'h10 ;
            rom[4402] = 8'hf6 ;
            rom[4403] = 8'h07 ;
            rom[4404] = 8'h03 ;
            rom[4405] = 8'he9 ;
            rom[4406] = 8'h0c ;
            rom[4407] = 8'h00 ;
            rom[4408] = 8'hf9 ;
            rom[4409] = 8'hdd ;
            rom[4410] = 8'h00 ;
            rom[4411] = 8'hf4 ;
            rom[4412] = 8'h09 ;
            rom[4413] = 8'h0c ;
            rom[4414] = 8'hf5 ;
            rom[4415] = 8'h0a ;
            rom[4416] = 8'h27 ;
            rom[4417] = 8'hf2 ;
            rom[4418] = 8'h07 ;
            rom[4419] = 8'hfb ;
            rom[4420] = 8'hed ;
            rom[4421] = 8'h04 ;
            rom[4422] = 8'h07 ;
            rom[4423] = 8'h01 ;
            rom[4424] = 8'h07 ;
            rom[4425] = 8'hf2 ;
            rom[4426] = 8'he9 ;
            rom[4427] = 8'h14 ;
            rom[4428] = 8'h0d ;
            rom[4429] = 8'hee ;
            rom[4430] = 8'hfc ;
            rom[4431] = 8'h21 ;
            rom[4432] = 8'h14 ;
            rom[4433] = 8'h00 ;
            rom[4434] = 8'hea ;
            rom[4435] = 8'h06 ;
            rom[4436] = 8'h0b ;
            rom[4437] = 8'h20 ;
            rom[4438] = 8'h21 ;
            rom[4439] = 8'hf8 ;
            rom[4440] = 8'hdf ;
            rom[4441] = 8'h15 ;
            rom[4442] = 8'hee ;
            rom[4443] = 8'h00 ;
            rom[4444] = 8'h0a ;
            rom[4445] = 8'h01 ;
            rom[4446] = 8'he6 ;
            rom[4447] = 8'hf4 ;
            rom[4448] = 8'h06 ;
            rom[4449] = 8'h08 ;
            rom[4450] = 8'hb6 ;
            rom[4451] = 8'hf9 ;
            rom[4452] = 8'hd5 ;
            rom[4453] = 8'hf5 ;
            rom[4454] = 8'h0c ;
            rom[4455] = 8'h1e ;
            rom[4456] = 8'hf8 ;
            rom[4457] = 8'h08 ;
            rom[4458] = 8'h19 ;
            rom[4459] = 8'hb1 ;
            rom[4460] = 8'hfd ;
            rom[4461] = 8'hf8 ;
            rom[4462] = 8'hfa ;
            rom[4463] = 8'hf1 ;
            rom[4464] = 8'hfc ;
            rom[4465] = 8'heb ;
            rom[4466] = 8'hfa ;
            rom[4467] = 8'hf2 ;
            rom[4468] = 8'h18 ;
            rom[4469] = 8'h04 ;
            rom[4470] = 8'hdd ;
            rom[4471] = 8'hfc ;
            rom[4472] = 8'hf2 ;
            rom[4473] = 8'hf7 ;
            rom[4474] = 8'hef ;
            rom[4475] = 8'hf3 ;
            rom[4476] = 8'h0a ;
            rom[4477] = 8'hf5 ;
            rom[4478] = 8'h07 ;
            rom[4479] = 8'he4 ;
            rom[4480] = 8'hfb ;
            rom[4481] = 8'h16 ;
            rom[4482] = 8'h05 ;
            rom[4483] = 8'hfe ;
            rom[4484] = 8'h08 ;
            rom[4485] = 8'hfb ;
            rom[4486] = 8'hf1 ;
            rom[4487] = 8'h0e ;
            rom[4488] = 8'h00 ;
            rom[4489] = 8'h04 ;
            rom[4490] = 8'hec ;
            rom[4491] = 8'hef ;
            rom[4492] = 8'hf9 ;
            rom[4493] = 8'hf4 ;
            rom[4494] = 8'h03 ;
            rom[4495] = 8'he8 ;
            rom[4496] = 8'hff ;
            rom[4497] = 8'h01 ;
            rom[4498] = 8'h11 ;
            rom[4499] = 8'h09 ;
            rom[4500] = 8'h01 ;
            rom[4501] = 8'h05 ;
            rom[4502] = 8'h0e ;
            rom[4503] = 8'hf1 ;
            rom[4504] = 8'hfa ;
            rom[4505] = 8'hf3 ;
            rom[4506] = 8'h0c ;
            rom[4507] = 8'hfd ;
            rom[4508] = 8'hd3 ;
            rom[4509] = 8'h1c ;
            rom[4510] = 8'hf9 ;
            rom[4511] = 8'hd2 ;
            rom[4512] = 8'h1e ;
            rom[4513] = 8'h23 ;
            rom[4514] = 8'h00 ;
            rom[4515] = 8'hd2 ;
            rom[4516] = 8'hfb ;
            rom[4517] = 8'h06 ;
            rom[4518] = 8'h10 ;
            rom[4519] = 8'h0f ;
            rom[4520] = 8'h09 ;
            rom[4521] = 8'h11 ;
            rom[4522] = 8'h1c ;
            rom[4523] = 8'hfe ;
            rom[4524] = 8'h18 ;
            rom[4525] = 8'hd7 ;
            rom[4526] = 8'h02 ;
            rom[4527] = 8'hfc ;
            rom[4528] = 8'hf3 ;
            rom[4529] = 8'h1a ;
            rom[4530] = 8'hf1 ;
            rom[4531] = 8'h1b ;
            rom[4532] = 8'h0c ;
            rom[4533] = 8'h18 ;
            rom[4534] = 8'h0b ;
            rom[4535] = 8'h0f ;
            rom[4536] = 8'hf8 ;
            rom[4537] = 8'h16 ;
            rom[4538] = 8'hdb ;
            rom[4539] = 8'h11 ;
            rom[4540] = 8'he8 ;
            rom[4541] = 8'hf5 ;
            rom[4542] = 8'hef ;
            rom[4543] = 8'hd9 ;
            rom[4544] = 8'h0c ;
            rom[4545] = 8'h09 ;
            rom[4546] = 8'h0a ;
            rom[4547] = 8'hf8 ;
            rom[4548] = 8'hfd ;
            rom[4549] = 8'h09 ;
            rom[4550] = 8'he7 ;
            rom[4551] = 8'h0b ;
            rom[4552] = 8'h35 ;
            rom[4553] = 8'h05 ;
            rom[4554] = 8'hf2 ;
            rom[4555] = 8'h07 ;
            rom[4556] = 8'h12 ;
            rom[4557] = 8'hf6 ;
            rom[4558] = 8'hec ;
            rom[4559] = 8'hf0 ;
            rom[4560] = 8'hf7 ;
            rom[4561] = 8'hfb ;
            rom[4562] = 8'he8 ;
            rom[4563] = 8'hfd ;
            rom[4564] = 8'h06 ;
            rom[4565] = 8'hcf ;
            rom[4566] = 8'h29 ;
            rom[4567] = 8'hcc ;
            rom[4568] = 8'h03 ;
            rom[4569] = 8'h00 ;
            rom[4570] = 8'h18 ;
            rom[4571] = 8'h08 ;
            rom[4572] = 8'he6 ;
            rom[4573] = 8'h0e ;
            rom[4574] = 8'h08 ;
            rom[4575] = 8'h07 ;
            rom[4576] = 8'h19 ;
            rom[4577] = 8'hf2 ;
            rom[4578] = 8'h0d ;
            rom[4579] = 8'h0c ;
            rom[4580] = 8'hfb ;
            rom[4581] = 8'h0d ;
            rom[4582] = 8'hff ;
            rom[4583] = 8'h0b ;
            rom[4584] = 8'hfa ;
            rom[4585] = 8'h04 ;
            rom[4586] = 8'hef ;
            rom[4587] = 8'h12 ;
            rom[4588] = 8'h10 ;
            rom[4589] = 8'h08 ;
            rom[4590] = 8'hfc ;
            rom[4591] = 8'h11 ;
            rom[4592] = 8'hfd ;
            rom[4593] = 8'hf2 ;
            rom[4594] = 8'hf1 ;
            rom[4595] = 8'h10 ;
            rom[4596] = 8'hfc ;
            rom[4597] = 8'hea ;
            rom[4598] = 8'hdc ;
            rom[4599] = 8'hdd ;
            rom[4600] = 8'h21 ;
            rom[4601] = 8'h0a ;
            rom[4602] = 8'hcc ;
            rom[4603] = 8'hfe ;
            rom[4604] = 8'h10 ;
            rom[4605] = 8'hf9 ;
            rom[4606] = 8'h0d ;
            rom[4607] = 8'hdc ;
            rom[4608] = 8'hff ;
            rom[4609] = 8'he3 ;
            rom[4610] = 8'hf0 ;
            rom[4611] = 8'hf5 ;
            rom[4612] = 8'h0b ;
            rom[4613] = 8'h14 ;
            rom[4614] = 8'h04 ;
            rom[4615] = 8'hfa ;
            rom[4616] = 8'h0e ;
            rom[4617] = 8'h0d ;
            rom[4618] = 8'he5 ;
            rom[4619] = 8'hef ;
            rom[4620] = 8'h0a ;
            rom[4621] = 8'hf9 ;
            rom[4622] = 8'h19 ;
            rom[4623] = 8'h29 ;
            rom[4624] = 8'h1f ;
            rom[4625] = 8'h04 ;
            rom[4626] = 8'h08 ;
            rom[4627] = 8'heb ;
            rom[4628] = 8'hea ;
            rom[4629] = 8'hd1 ;
            rom[4630] = 8'h06 ;
            rom[4631] = 8'hff ;
            rom[4632] = 8'hf3 ;
            rom[4633] = 8'h23 ;
            rom[4634] = 8'h07 ;
            rom[4635] = 8'h11 ;
            rom[4636] = 8'h08 ;
            rom[4637] = 8'hf2 ;
            rom[4638] = 8'h00 ;
            rom[4639] = 8'hfd ;
            rom[4640] = 8'h03 ;
            rom[4641] = 8'h17 ;
            rom[4642] = 8'h10 ;
            rom[4643] = 8'h1b ;
            rom[4644] = 8'h1c ;
            rom[4645] = 8'h06 ;
            rom[4646] = 8'h04 ;
            rom[4647] = 8'he9 ;
            rom[4648] = 8'h02 ;
            rom[4649] = 8'hf6 ;
            rom[4650] = 8'h12 ;
            rom[4651] = 8'hec ;
            rom[4652] = 8'h00 ;
            rom[4653] = 8'hef ;
            rom[4654] = 8'h07 ;
            rom[4655] = 8'hf1 ;
            rom[4656] = 8'h15 ;
            rom[4657] = 8'hfd ;
            rom[4658] = 8'hfa ;
            rom[4659] = 8'h1f ;
            rom[4660] = 8'h17 ;
            rom[4661] = 8'hfc ;
            rom[4662] = 8'h07 ;
            rom[4663] = 8'he2 ;
            rom[4664] = 8'hff ;
            rom[4665] = 8'hf1 ;
            rom[4666] = 8'h05 ;
            rom[4667] = 8'hfc ;
            rom[4668] = 8'h08 ;
            rom[4669] = 8'h20 ;
            rom[4670] = 8'h10 ;
            rom[4671] = 8'h1a ;
            rom[4672] = 8'hf4 ;
            rom[4673] = 8'hd8 ;
            rom[4674] = 8'hfd ;
            rom[4675] = 8'h04 ;
            rom[4676] = 8'h1c ;
            rom[4677] = 8'hf5 ;
            rom[4678] = 8'h0d ;
            rom[4679] = 8'hf0 ;
            rom[4680] = 8'h1f ;
            rom[4681] = 8'h0f ;
            rom[4682] = 8'h0f ;
            rom[4683] = 8'hf9 ;
            rom[4684] = 8'h15 ;
            rom[4685] = 8'hfd ;
            rom[4686] = 8'hf9 ;
            rom[4687] = 8'h16 ;
            rom[4688] = 8'h14 ;
            rom[4689] = 8'h01 ;
            rom[4690] = 8'h09 ;
            rom[4691] = 8'h03 ;
            rom[4692] = 8'hf3 ;
            rom[4693] = 8'hec ;
            rom[4694] = 8'h06 ;
            rom[4695] = 8'hfe ;
            rom[4696] = 8'h12 ;
            rom[4697] = 8'h1c ;
            rom[4698] = 8'hff ;
            rom[4699] = 8'h15 ;
            rom[4700] = 8'h1d ;
            rom[4701] = 8'h08 ;
            rom[4702] = 8'h1b ;
            rom[4703] = 8'hf0 ;
            rom[4704] = 8'hf7 ;
            rom[4705] = 8'h1b ;
            rom[4706] = 8'h19 ;
            rom[4707] = 8'hf5 ;
            rom[4708] = 8'h2e ;
            rom[4709] = 8'h11 ;
            rom[4710] = 8'hf3 ;
            rom[4711] = 8'he9 ;
            rom[4712] = 8'h00 ;
            rom[4713] = 8'h0a ;
            rom[4714] = 8'h05 ;
            rom[4715] = 8'h05 ;
            rom[4716] = 8'hfb ;
            rom[4717] = 8'he7 ;
            rom[4718] = 8'h10 ;
            rom[4719] = 8'hfb ;
            rom[4720] = 8'h04 ;
            rom[4721] = 8'h00 ;
            rom[4722] = 8'h00 ;
            rom[4723] = 8'h1d ;
            rom[4724] = 8'h08 ;
            rom[4725] = 8'hfb ;
            rom[4726] = 8'h02 ;
            rom[4727] = 8'he5 ;
            rom[4728] = 8'h08 ;
            rom[4729] = 8'hef ;
            rom[4730] = 8'hf0 ;
            rom[4731] = 8'h15 ;
            rom[4732] = 8'h07 ;
            rom[4733] = 8'h05 ;
            rom[4734] = 8'h03 ;
            rom[4735] = 8'h1a ;
            rom[4736] = 8'hf1 ;
            rom[4737] = 8'hd1 ;
            rom[4738] = 8'hfa ;
            rom[4739] = 8'h04 ;
            rom[4740] = 8'hfe ;
            rom[4741] = 8'h1a ;
            rom[4742] = 8'h06 ;
            rom[4743] = 8'hdb ;
            rom[4744] = 8'h0f ;
            rom[4745] = 8'hfe ;
            rom[4746] = 8'hf5 ;
            rom[4747] = 8'heb ;
            rom[4748] = 8'hde ;
            rom[4749] = 8'h04 ;
            rom[4750] = 8'h0d ;
            rom[4751] = 8'h35 ;
            rom[4752] = 8'h07 ;
            rom[4753] = 8'hfd ;
            rom[4754] = 8'hfa ;
            rom[4755] = 8'h1c ;
            rom[4756] = 8'h05 ;
            rom[4757] = 8'hfa ;
            rom[4758] = 8'h1e ;
            rom[4759] = 8'hfa ;
            rom[4760] = 8'hf3 ;
            rom[4761] = 8'h02 ;
            rom[4762] = 8'h10 ;
            rom[4763] = 8'he0 ;
            rom[4764] = 8'h06 ;
            rom[4765] = 8'hec ;
            rom[4766] = 8'hfa ;
            rom[4767] = 8'he9 ;
            rom[4768] = 8'hf2 ;
            rom[4769] = 8'h10 ;
            rom[4770] = 8'h07 ;
            rom[4771] = 8'hfc ;
            rom[4772] = 8'hf3 ;
            rom[4773] = 8'hf9 ;
            rom[4774] = 8'hf2 ;
            rom[4775] = 8'h1b ;
            rom[4776] = 8'he1 ;
            rom[4777] = 8'h05 ;
            rom[4778] = 8'h1b ;
            rom[4779] = 8'h03 ;
            rom[4780] = 8'h18 ;
            rom[4781] = 8'h01 ;
            rom[4782] = 8'hf5 ;
            rom[4783] = 8'h05 ;
            rom[4784] = 8'he8 ;
            rom[4785] = 8'hf6 ;
            rom[4786] = 8'hf1 ;
            rom[4787] = 8'h10 ;
            rom[4788] = 8'h10 ;
            rom[4789] = 8'h00 ;
            rom[4790] = 8'he9 ;
            rom[4791] = 8'hcc ;
            rom[4792] = 8'hfc ;
            rom[4793] = 8'h17 ;
            rom[4794] = 8'h09 ;
            rom[4795] = 8'h05 ;
            rom[4796] = 8'h22 ;
            rom[4797] = 8'h04 ;
            rom[4798] = 8'hfc ;
            rom[4799] = 8'hee ;
            rom[4800] = 8'h01 ;
            rom[4801] = 8'h0f ;
            rom[4802] = 8'heb ;
            rom[4803] = 8'heb ;
            rom[4804] = 8'hf8 ;
            rom[4805] = 8'h15 ;
            rom[4806] = 8'h18 ;
            rom[4807] = 8'h1f ;
            rom[4808] = 8'h22 ;
            rom[4809] = 8'h03 ;
            rom[4810] = 8'hf2 ;
            rom[4811] = 8'hf9 ;
            rom[4812] = 8'h1c ;
            rom[4813] = 8'hec ;
            rom[4814] = 8'h2b ;
            rom[4815] = 8'h20 ;
            rom[4816] = 8'h24 ;
            rom[4817] = 8'hfb ;
            rom[4818] = 8'hf9 ;
            rom[4819] = 8'h07 ;
            rom[4820] = 8'hf8 ;
            rom[4821] = 8'h16 ;
            rom[4822] = 8'h0c ;
            rom[4823] = 8'hf9 ;
            rom[4824] = 8'hf9 ;
            rom[4825] = 8'h03 ;
            rom[4826] = 8'h07 ;
            rom[4827] = 8'hfe ;
            rom[4828] = 8'h04 ;
            rom[4829] = 8'hcb ;
            rom[4830] = 8'h0d ;
            rom[4831] = 8'hf6 ;
            rom[4832] = 8'hea ;
            rom[4833] = 8'h27 ;
            rom[4834] = 8'h26 ;
            rom[4835] = 8'hf4 ;
            rom[4836] = 8'hdc ;
            rom[4837] = 8'hfd ;
            rom[4838] = 8'h11 ;
            rom[4839] = 8'hf4 ;
            rom[4840] = 8'hd7 ;
            rom[4841] = 8'h19 ;
            rom[4842] = 8'hd8 ;
            rom[4843] = 8'hee ;
            rom[4844] = 8'hee ;
            rom[4845] = 8'he4 ;
            rom[4846] = 8'h0c ;
            rom[4847] = 8'h15 ;
            rom[4848] = 8'he9 ;
            rom[4849] = 8'hfe ;
            rom[4850] = 8'h1e ;
            rom[4851] = 8'he9 ;
            rom[4852] = 8'hfc ;
            rom[4853] = 8'hfc ;
            rom[4854] = 8'hf1 ;
            rom[4855] = 8'hfd ;
            rom[4856] = 8'hdc ;
            rom[4857] = 8'h0c ;
            rom[4858] = 8'hf9 ;
            rom[4859] = 8'hf5 ;
            rom[4860] = 8'h01 ;
            rom[4861] = 8'h01 ;
            rom[4862] = 8'hf1 ;
            rom[4863] = 8'h0a ;
            rom[4864] = 8'h00 ;
            rom[4865] = 8'h12 ;
            rom[4866] = 8'h09 ;
            rom[4867] = 8'h02 ;
            rom[4868] = 8'h03 ;
            rom[4869] = 8'h04 ;
            rom[4870] = 8'hd7 ;
            rom[4871] = 8'h0d ;
            rom[4872] = 8'h12 ;
            rom[4873] = 8'h0b ;
            rom[4874] = 8'hef ;
            rom[4875] = 8'hff ;
            rom[4876] = 8'h07 ;
            rom[4877] = 8'hea ;
            rom[4878] = 8'hec ;
            rom[4879] = 8'h07 ;
            rom[4880] = 8'h03 ;
            rom[4881] = 8'hfa ;
            rom[4882] = 8'h1b ;
            rom[4883] = 8'he7 ;
            rom[4884] = 8'he4 ;
            rom[4885] = 8'h05 ;
            rom[4886] = 8'h19 ;
            rom[4887] = 8'hf6 ;
            rom[4888] = 8'he2 ;
            rom[4889] = 8'h07 ;
            rom[4890] = 8'h14 ;
            rom[4891] = 8'he7 ;
            rom[4892] = 8'hf1 ;
            rom[4893] = 8'h15 ;
            rom[4894] = 8'hfe ;
            rom[4895] = 8'hfd ;
            rom[4896] = 8'h11 ;
            rom[4897] = 8'h06 ;
            rom[4898] = 8'h0f ;
            rom[4899] = 8'h1b ;
            rom[4900] = 8'hdc ;
            rom[4901] = 8'h0b ;
            rom[4902] = 8'hff ;
            rom[4903] = 8'h19 ;
            rom[4904] = 8'h0c ;
            rom[4905] = 8'hf4 ;
            rom[4906] = 8'h0f ;
            rom[4907] = 8'h21 ;
            rom[4908] = 8'hff ;
            rom[4909] = 8'hc2 ;
            rom[4910] = 8'h10 ;
            rom[4911] = 8'h11 ;
            rom[4912] = 8'he9 ;
            rom[4913] = 8'h0c ;
            rom[4914] = 8'hf6 ;
            rom[4915] = 8'h0b ;
            rom[4916] = 8'h04 ;
            rom[4917] = 8'he8 ;
            rom[4918] = 8'h16 ;
            rom[4919] = 8'hfd ;
            rom[4920] = 8'h0e ;
            rom[4921] = 8'h0f ;
            rom[4922] = 8'hca ;
            rom[4923] = 8'h16 ;
            rom[4924] = 8'hed ;
            rom[4925] = 8'hf9 ;
            rom[4926] = 8'he3 ;
            rom[4927] = 8'hd2 ;
            rom[4928] = 8'hfa ;
            rom[4929] = 8'h14 ;
            rom[4930] = 8'hed ;
            rom[4931] = 8'hf9 ;
            rom[4932] = 8'he5 ;
            rom[4933] = 8'hfc ;
            rom[4934] = 8'h1d ;
            rom[4935] = 8'hfc ;
            rom[4936] = 8'hfe ;
            rom[4937] = 8'h09 ;
            rom[4938] = 8'hf1 ;
            rom[4939] = 8'hea ;
            rom[4940] = 8'hd6 ;
            rom[4941] = 8'hf2 ;
            rom[4942] = 8'h0b ;
            rom[4943] = 8'h14 ;
            rom[4944] = 8'hfd ;
            rom[4945] = 8'h02 ;
            rom[4946] = 8'h17 ;
            rom[4947] = 8'hca ;
            rom[4948] = 8'hfa ;
            rom[4949] = 8'hf0 ;
            rom[4950] = 8'h23 ;
            rom[4951] = 8'h1e ;
            rom[4952] = 8'h25 ;
            rom[4953] = 8'h0d ;
            rom[4954] = 8'h13 ;
            rom[4955] = 8'hf9 ;
            rom[4956] = 8'hee ;
            rom[4957] = 8'hfd ;
            rom[4958] = 8'hfd ;
            rom[4959] = 8'hf7 ;
            rom[4960] = 8'he3 ;
            rom[4961] = 8'he6 ;
            rom[4962] = 8'hf2 ;
            rom[4963] = 8'h12 ;
            rom[4964] = 8'h06 ;
            rom[4965] = 8'hf7 ;
            rom[4966] = 8'h09 ;
            rom[4967] = 8'he1 ;
            rom[4968] = 8'he7 ;
            rom[4969] = 8'h1b ;
            rom[4970] = 8'h01 ;
            rom[4971] = 8'he9 ;
            rom[4972] = 8'hfc ;
            rom[4973] = 8'he7 ;
            rom[4974] = 8'h14 ;
            rom[4975] = 8'hf8 ;
            rom[4976] = 8'h1d ;
            rom[4977] = 8'h03 ;
            rom[4978] = 8'h11 ;
            rom[4979] = 8'hf6 ;
            rom[4980] = 8'h1c ;
            rom[4981] = 8'hfe ;
            rom[4982] = 8'hfb ;
            rom[4983] = 8'he8 ;
            rom[4984] = 8'hf1 ;
            rom[4985] = 8'hf9 ;
            rom[4986] = 8'hef ;
            rom[4987] = 8'h11 ;
            rom[4988] = 8'hee ;
            rom[4989] = 8'he2 ;
            rom[4990] = 8'hee ;
            rom[4991] = 8'hfb ;
            rom[4992] = 8'h08 ;
            rom[4993] = 8'h0e ;
            rom[4994] = 8'h08 ;
            rom[4995] = 8'h0c ;
            rom[4996] = 8'hf8 ;
            rom[4997] = 8'hd8 ;
            rom[4998] = 8'h0c ;
            rom[4999] = 8'hfd ;
            rom[5000] = 8'h2d ;
            rom[5001] = 8'h0d ;
            rom[5002] = 8'hff ;
            rom[5003] = 8'hf1 ;
            rom[5004] = 8'hec ;
            rom[5005] = 8'he7 ;
            rom[5006] = 8'h0c ;
            rom[5007] = 8'hf7 ;
            rom[5008] = 8'hf7 ;
            rom[5009] = 8'hf9 ;
            rom[5010] = 8'hf5 ;
            rom[5011] = 8'hfa ;
            rom[5012] = 8'h02 ;
            rom[5013] = 8'hf1 ;
            rom[5014] = 8'h0e ;
            rom[5015] = 8'h22 ;
            rom[5016] = 8'hfd ;
            rom[5017] = 8'h0e ;
            rom[5018] = 8'h00 ;
            rom[5019] = 8'h2a ;
            rom[5020] = 8'h12 ;
            rom[5021] = 8'h16 ;
            rom[5022] = 8'h02 ;
            rom[5023] = 8'hfa ;
            rom[5024] = 8'hfd ;
            rom[5025] = 8'h17 ;
            rom[5026] = 8'h09 ;
            rom[5027] = 8'h04 ;
            rom[5028] = 8'hff ;
            rom[5029] = 8'he7 ;
            rom[5030] = 8'hf2 ;
            rom[5031] = 8'he9 ;
            rom[5032] = 8'hff ;
            rom[5033] = 8'h07 ;
            rom[5034] = 8'heb ;
            rom[5035] = 8'hfc ;
            rom[5036] = 8'he3 ;
            rom[5037] = 8'hd9 ;
            rom[5038] = 8'hf1 ;
            rom[5039] = 8'he6 ;
            rom[5040] = 8'h13 ;
            rom[5041] = 8'hf1 ;
            rom[5042] = 8'h20 ;
            rom[5043] = 8'he7 ;
            rom[5044] = 8'he8 ;
            rom[5045] = 8'hf7 ;
            rom[5046] = 8'h08 ;
            rom[5047] = 8'h10 ;
            rom[5048] = 8'h03 ;
            rom[5049] = 8'h13 ;
            rom[5050] = 8'hff ;
            rom[5051] = 8'he0 ;
            rom[5052] = 8'h0f ;
            rom[5053] = 8'hfc ;
            rom[5054] = 8'he6 ;
            rom[5055] = 8'hf5 ;
            rom[5056] = 8'h07 ;
            rom[5057] = 8'h03 ;
            rom[5058] = 8'h06 ;
            rom[5059] = 8'h11 ;
            rom[5060] = 8'he1 ;
            rom[5061] = 8'h03 ;
            rom[5062] = 8'h00 ;
            rom[5063] = 8'h01 ;
            rom[5064] = 8'h10 ;
            rom[5065] = 8'h04 ;
            rom[5066] = 8'hf9 ;
            rom[5067] = 8'hdb ;
            rom[5068] = 8'h00 ;
            rom[5069] = 8'h00 ;
            rom[5070] = 8'h0c ;
            rom[5071] = 8'h0e ;
            rom[5072] = 8'h0a ;
            rom[5073] = 8'hc7 ;
            rom[5074] = 8'hf8 ;
            rom[5075] = 8'hda ;
            rom[5076] = 8'hf7 ;
            rom[5077] = 8'hed ;
            rom[5078] = 8'h0f ;
            rom[5079] = 8'hfe ;
            rom[5080] = 8'hf9 ;
            rom[5081] = 8'hf5 ;
            rom[5082] = 8'h08 ;
            rom[5083] = 8'h0d ;
            rom[5084] = 8'h00 ;
            rom[5085] = 8'h0a ;
            rom[5086] = 8'h15 ;
            rom[5087] = 8'hfd ;
            rom[5088] = 8'hf7 ;
            rom[5089] = 8'h30 ;
            rom[5090] = 8'h1f ;
            rom[5091] = 8'hfd ;
            rom[5092] = 8'hf9 ;
            rom[5093] = 8'h01 ;
            rom[5094] = 8'hf4 ;
            rom[5095] = 8'h00 ;
            rom[5096] = 8'hff ;
            rom[5097] = 8'hff ;
            rom[5098] = 8'he4 ;
            rom[5099] = 8'h1b ;
            rom[5100] = 8'hc4 ;
            rom[5101] = 8'hc9 ;
            rom[5102] = 8'h19 ;
            rom[5103] = 8'h18 ;
            rom[5104] = 8'he4 ;
            rom[5105] = 8'hff ;
            rom[5106] = 8'h20 ;
            rom[5107] = 8'hfa ;
            rom[5108] = 8'h06 ;
            rom[5109] = 8'he0 ;
            rom[5110] = 8'h01 ;
            rom[5111] = 8'hea ;
            rom[5112] = 8'h16 ;
            rom[5113] = 8'h0c ;
            rom[5114] = 8'hef ;
            rom[5115] = 8'hf7 ;
            rom[5116] = 8'hf4 ;
            rom[5117] = 8'h1a ;
            rom[5118] = 8'he3 ;
            rom[5119] = 8'h04 ;
            rom[5120] = 8'h07 ;
            rom[5121] = 8'h0c ;
            rom[5122] = 8'h0b ;
            rom[5123] = 8'h18 ;
            rom[5124] = 8'h0e ;
            rom[5125] = 8'hdb ;
            rom[5126] = 8'hc0 ;
            rom[5127] = 8'hea ;
            rom[5128] = 8'hf5 ;
            rom[5129] = 8'h0b ;
            rom[5130] = 8'h08 ;
            rom[5131] = 8'h09 ;
            rom[5132] = 8'h06 ;
            rom[5133] = 8'he0 ;
            rom[5134] = 8'he8 ;
            rom[5135] = 8'h14 ;
            rom[5136] = 8'hf8 ;
            rom[5137] = 8'hff ;
            rom[5138] = 8'hfe ;
            rom[5139] = 8'hfa ;
            rom[5140] = 8'h03 ;
            rom[5141] = 8'h23 ;
            rom[5142] = 8'hf4 ;
            rom[5143] = 8'h00 ;
            rom[5144] = 8'hfe ;
            rom[5145] = 8'h1b ;
            rom[5146] = 8'he9 ;
            rom[5147] = 8'he0 ;
            rom[5148] = 8'hed ;
            rom[5149] = 8'h1c ;
            rom[5150] = 8'he9 ;
            rom[5151] = 8'hf6 ;
            rom[5152] = 8'h33 ;
            rom[5153] = 8'h0a ;
            rom[5154] = 8'h0d ;
            rom[5155] = 8'he3 ;
            rom[5156] = 8'hf9 ;
            rom[5157] = 8'hf9 ;
            rom[5158] = 8'h17 ;
            rom[5159] = 8'hf3 ;
            rom[5160] = 8'h0a ;
            rom[5161] = 8'h0c ;
            rom[5162] = 8'hf9 ;
            rom[5163] = 8'h08 ;
            rom[5164] = 8'hfb ;
            rom[5165] = 8'h08 ;
            rom[5166] = 8'h22 ;
            rom[5167] = 8'h0e ;
            rom[5168] = 8'he9 ;
            rom[5169] = 8'h09 ;
            rom[5170] = 8'hfe ;
            rom[5171] = 8'h17 ;
            rom[5172] = 8'h05 ;
            rom[5173] = 8'hd4 ;
            rom[5174] = 8'h03 ;
            rom[5175] = 8'h1a ;
            rom[5176] = 8'hf2 ;
            rom[5177] = 8'hf4 ;
            rom[5178] = 8'heb ;
            rom[5179] = 8'hfa ;
            rom[5180] = 8'h0b ;
            rom[5181] = 8'hf0 ;
            rom[5182] = 8'hff ;
            rom[5183] = 8'hf8 ;
            rom[5184] = 8'hea ;
            rom[5185] = 8'h02 ;
            rom[5186] = 8'hf2 ;
            rom[5187] = 8'hff ;
            rom[5188] = 8'h0c ;
            rom[5189] = 8'h19 ;
            rom[5190] = 8'h07 ;
            rom[5191] = 8'h12 ;
            rom[5192] = 8'h24 ;
            rom[5193] = 8'h0a ;
            rom[5194] = 8'heb ;
            rom[5195] = 8'h0b ;
            rom[5196] = 8'h07 ;
            rom[5197] = 8'h15 ;
            rom[5198] = 8'hf5 ;
            rom[5199] = 8'he8 ;
            rom[5200] = 8'hf0 ;
            rom[5201] = 8'hf6 ;
            rom[5202] = 8'hf0 ;
            rom[5203] = 8'h07 ;
            rom[5204] = 8'hfe ;
            rom[5205] = 8'h06 ;
            rom[5206] = 8'h0a ;
            rom[5207] = 8'h11 ;
            rom[5208] = 8'hfe ;
            rom[5209] = 8'h15 ;
            rom[5210] = 8'h0e ;
            rom[5211] = 8'h10 ;
            rom[5212] = 8'hfe ;
            rom[5213] = 8'hfc ;
            rom[5214] = 8'h12 ;
            rom[5215] = 8'h09 ;
            rom[5216] = 8'h22 ;
            rom[5217] = 8'hed ;
            rom[5218] = 8'h0f ;
            rom[5219] = 8'h17 ;
            rom[5220] = 8'h0b ;
            rom[5221] = 8'he3 ;
            rom[5222] = 8'hff ;
            rom[5223] = 8'hf9 ;
            rom[5224] = 8'hee ;
            rom[5225] = 8'hea ;
            rom[5226] = 8'h00 ;
            rom[5227] = 8'hfc ;
            rom[5228] = 8'h02 ;
            rom[5229] = 8'h06 ;
            rom[5230] = 8'h04 ;
            rom[5231] = 8'h0b ;
            rom[5232] = 8'hfa ;
            rom[5233] = 8'h0e ;
            rom[5234] = 8'hde ;
            rom[5235] = 8'h1e ;
            rom[5236] = 8'hf4 ;
            rom[5237] = 8'hea ;
            rom[5238] = 8'h08 ;
            rom[5239] = 8'he9 ;
            rom[5240] = 8'hd4 ;
            rom[5241] = 8'he4 ;
            rom[5242] = 8'hfa ;
            rom[5243] = 8'hf6 ;
            rom[5244] = 8'h1e ;
            rom[5245] = 8'h19 ;
            rom[5246] = 8'h0e ;
            rom[5247] = 8'hf2 ;
            rom[5248] = 8'he7 ;
            rom[5249] = 8'hfd ;
            rom[5250] = 8'hf6 ;
            rom[5251] = 8'h1a ;
            rom[5252] = 8'h06 ;
            rom[5253] = 8'hfc ;
            rom[5254] = 8'h1b ;
            rom[5255] = 8'hff ;
            rom[5256] = 8'h0d ;
            rom[5257] = 8'h1d ;
            rom[5258] = 8'hfc ;
            rom[5259] = 8'h03 ;
            rom[5260] = 8'hfe ;
            rom[5261] = 8'he8 ;
            rom[5262] = 8'hfd ;
            rom[5263] = 8'hfd ;
            rom[5264] = 8'hf6 ;
            rom[5265] = 8'h02 ;
            rom[5266] = 8'hf9 ;
            rom[5267] = 8'h05 ;
            rom[5268] = 8'hfd ;
            rom[5269] = 8'h01 ;
            rom[5270] = 8'h0b ;
            rom[5271] = 8'h26 ;
            rom[5272] = 8'h08 ;
            rom[5273] = 8'h00 ;
            rom[5274] = 8'h02 ;
            rom[5275] = 8'hf2 ;
            rom[5276] = 8'hf1 ;
            rom[5277] = 8'h17 ;
            rom[5278] = 8'h0d ;
            rom[5279] = 8'hd8 ;
            rom[5280] = 8'h08 ;
            rom[5281] = 8'hef ;
            rom[5282] = 8'hee ;
            rom[5283] = 8'h16 ;
            rom[5284] = 8'he5 ;
            rom[5285] = 8'h00 ;
            rom[5286] = 8'h09 ;
            rom[5287] = 8'hfd ;
            rom[5288] = 8'h0e ;
            rom[5289] = 8'hf8 ;
            rom[5290] = 8'h1a ;
            rom[5291] = 8'h05 ;
            rom[5292] = 8'h19 ;
            rom[5293] = 8'h14 ;
            rom[5294] = 8'h13 ;
            rom[5295] = 8'hef ;
            rom[5296] = 8'hfb ;
            rom[5297] = 8'h0e ;
            rom[5298] = 8'h06 ;
            rom[5299] = 8'hff ;
            rom[5300] = 8'hf0 ;
            rom[5301] = 8'h0d ;
            rom[5302] = 8'h16 ;
            rom[5303] = 8'h04 ;
            rom[5304] = 8'h01 ;
            rom[5305] = 8'h05 ;
            rom[5306] = 8'h01 ;
            rom[5307] = 8'hfa ;
            rom[5308] = 8'hef ;
            rom[5309] = 8'h22 ;
            rom[5310] = 8'hf2 ;
            rom[5311] = 8'hcf ;
            rom[5312] = 8'he8 ;
            rom[5313] = 8'h11 ;
            rom[5314] = 8'he7 ;
            rom[5315] = 8'hfe ;
            rom[5316] = 8'h07 ;
            rom[5317] = 8'h0b ;
            rom[5318] = 8'h03 ;
            rom[5319] = 8'h03 ;
            rom[5320] = 8'h05 ;
            rom[5321] = 8'hf7 ;
            rom[5322] = 8'ha5 ;
            rom[5323] = 8'hf6 ;
            rom[5324] = 8'hde ;
            rom[5325] = 8'h05 ;
            rom[5326] = 8'hef ;
            rom[5327] = 8'h26 ;
            rom[5328] = 8'h24 ;
            rom[5329] = 8'hf5 ;
            rom[5330] = 8'h08 ;
            rom[5331] = 8'hec ;
            rom[5332] = 8'hf7 ;
            rom[5333] = 8'h0d ;
            rom[5334] = 8'hfb ;
            rom[5335] = 8'h02 ;
            rom[5336] = 8'h06 ;
            rom[5337] = 8'h02 ;
            rom[5338] = 8'h22 ;
            rom[5339] = 8'h14 ;
            rom[5340] = 8'h02 ;
            rom[5341] = 8'he5 ;
            rom[5342] = 8'h1d ;
            rom[5343] = 8'he9 ;
            rom[5344] = 8'hf8 ;
            rom[5345] = 8'h0d ;
            rom[5346] = 8'h24 ;
            rom[5347] = 8'h1a ;
            rom[5348] = 8'he9 ;
            rom[5349] = 8'h04 ;
            rom[5350] = 8'he1 ;
            rom[5351] = 8'h08 ;
            rom[5352] = 8'h1b ;
            rom[5353] = 8'h03 ;
            rom[5354] = 8'he1 ;
            rom[5355] = 8'he9 ;
            rom[5356] = 8'h04 ;
            rom[5357] = 8'hf6 ;
            rom[5358] = 8'hdc ;
            rom[5359] = 8'hfa ;
            rom[5360] = 8'h0c ;
            rom[5361] = 8'hf2 ;
            rom[5362] = 8'he2 ;
            rom[5363] = 8'hf9 ;
            rom[5364] = 8'h0a ;
            rom[5365] = 8'h11 ;
            rom[5366] = 8'hf6 ;
            rom[5367] = 8'h0a ;
            rom[5368] = 8'hd9 ;
            rom[5369] = 8'h21 ;
            rom[5370] = 8'hd9 ;
            rom[5371] = 8'hed ;
            rom[5372] = 8'h06 ;
            rom[5373] = 8'h0c ;
            rom[5374] = 8'hfc ;
            rom[5375] = 8'h06 ;
            rom[5376] = 8'h0c ;
            rom[5377] = 8'he6 ;
            rom[5378] = 8'h00 ;
            rom[5379] = 8'h11 ;
            rom[5380] = 8'h0b ;
            rom[5381] = 8'hd3 ;
            rom[5382] = 8'hfa ;
            rom[5383] = 8'he3 ;
            rom[5384] = 8'h0a ;
            rom[5385] = 8'h11 ;
            rom[5386] = 8'h0e ;
            rom[5387] = 8'h0c ;
            rom[5388] = 8'h32 ;
            rom[5389] = 8'he9 ;
            rom[5390] = 8'hfd ;
            rom[5391] = 8'h0f ;
            rom[5392] = 8'h08 ;
            rom[5393] = 8'h24 ;
            rom[5394] = 8'hef ;
            rom[5395] = 8'h02 ;
            rom[5396] = 8'he7 ;
            rom[5397] = 8'h21 ;
            rom[5398] = 8'hf9 ;
            rom[5399] = 8'hf3 ;
            rom[5400] = 8'h16 ;
            rom[5401] = 8'h13 ;
            rom[5402] = 8'he5 ;
            rom[5403] = 8'he9 ;
            rom[5404] = 8'h15 ;
            rom[5405] = 8'h0e ;
            rom[5406] = 8'he7 ;
            rom[5407] = 8'hf3 ;
            rom[5408] = 8'h11 ;
            rom[5409] = 8'hf3 ;
            rom[5410] = 8'hf3 ;
            rom[5411] = 8'hea ;
            rom[5412] = 8'h09 ;
            rom[5413] = 8'hfb ;
            rom[5414] = 8'h1e ;
            rom[5415] = 8'hee ;
            rom[5416] = 8'h10 ;
            rom[5417] = 8'he9 ;
            rom[5418] = 8'hfa ;
            rom[5419] = 8'h03 ;
            rom[5420] = 8'h04 ;
            rom[5421] = 8'hf0 ;
            rom[5422] = 8'h19 ;
            rom[5423] = 8'hf0 ;
            rom[5424] = 8'h20 ;
            rom[5425] = 8'hf6 ;
            rom[5426] = 8'hff ;
            rom[5427] = 8'h24 ;
            rom[5428] = 8'h0b ;
            rom[5429] = 8'h0a ;
            rom[5430] = 8'hfb ;
            rom[5431] = 8'hfc ;
            rom[5432] = 8'hfe ;
            rom[5433] = 8'hcf ;
            rom[5434] = 8'h0c ;
            rom[5435] = 8'h07 ;
            rom[5436] = 8'h23 ;
            rom[5437] = 8'h14 ;
            rom[5438] = 8'he2 ;
            rom[5439] = 8'h1b ;
            rom[5440] = 8'h16 ;
            rom[5441] = 8'hd4 ;
            rom[5442] = 8'h1c ;
            rom[5443] = 8'h0e ;
            rom[5444] = 8'h02 ;
            rom[5445] = 8'he0 ;
            rom[5446] = 8'hf7 ;
            rom[5447] = 8'h0d ;
            rom[5448] = 8'h0e ;
            rom[5449] = 8'hf1 ;
            rom[5450] = 8'hef ;
            rom[5451] = 8'hf0 ;
            rom[5452] = 8'h03 ;
            rom[5453] = 8'h1a ;
            rom[5454] = 8'hfe ;
            rom[5455] = 8'h01 ;
            rom[5456] = 8'h0c ;
            rom[5457] = 8'hed ;
            rom[5458] = 8'hdd ;
            rom[5459] = 8'h10 ;
            rom[5460] = 8'h01 ;
            rom[5461] = 8'h09 ;
            rom[5462] = 8'h0e ;
            rom[5463] = 8'h20 ;
            rom[5464] = 8'h1b ;
            rom[5465] = 8'hfb ;
            rom[5466] = 8'h24 ;
            rom[5467] = 8'h08 ;
            rom[5468] = 8'h1a ;
            rom[5469] = 8'hdb ;
            rom[5470] = 8'he7 ;
            rom[5471] = 8'h09 ;
            rom[5472] = 8'h2a ;
            rom[5473] = 8'h09 ;
            rom[5474] = 8'h04 ;
            rom[5475] = 8'h11 ;
            rom[5476] = 8'hc4 ;
            rom[5477] = 8'h1b ;
            rom[5478] = 8'h15 ;
            rom[5479] = 8'hed ;
            rom[5480] = 8'hed ;
            rom[5481] = 8'h26 ;
            rom[5482] = 8'h0d ;
            rom[5483] = 8'he5 ;
            rom[5484] = 8'h16 ;
            rom[5485] = 8'h0d ;
            rom[5486] = 8'h0d ;
            rom[5487] = 8'h15 ;
            rom[5488] = 8'h05 ;
            rom[5489] = 8'hfc ;
            rom[5490] = 8'h23 ;
            rom[5491] = 8'h0b ;
            rom[5492] = 8'h04 ;
            rom[5493] = 8'hf6 ;
            rom[5494] = 8'h0e ;
            rom[5495] = 8'h07 ;
            rom[5496] = 8'h00 ;
            rom[5497] = 8'h00 ;
            rom[5498] = 8'h12 ;
            rom[5499] = 8'hc6 ;
            rom[5500] = 8'h1e ;
            rom[5501] = 8'hf1 ;
            rom[5502] = 8'h0f ;
            rom[5503] = 8'hfd ;
            rom[5504] = 8'hf4 ;
            rom[5505] = 8'hd3 ;
            rom[5506] = 8'hf6 ;
            rom[5507] = 8'he8 ;
            rom[5508] = 8'hf8 ;
            rom[5509] = 8'h16 ;
            rom[5510] = 8'h03 ;
            rom[5511] = 8'hea ;
            rom[5512] = 8'h0a ;
            rom[5513] = 8'hfc ;
            rom[5514] = 8'heb ;
            rom[5515] = 8'h02 ;
            rom[5516] = 8'hfa ;
            rom[5517] = 8'hf2 ;
            rom[5518] = 8'he6 ;
            rom[5519] = 8'h21 ;
            rom[5520] = 8'h0c ;
            rom[5521] = 8'hfd ;
            rom[5522] = 8'hf0 ;
            rom[5523] = 8'hdb ;
            rom[5524] = 8'hf9 ;
            rom[5525] = 8'hf4 ;
            rom[5526] = 8'h1b ;
            rom[5527] = 8'hea ;
            rom[5528] = 8'hdf ;
            rom[5529] = 8'h0b ;
            rom[5530] = 8'h0f ;
            rom[5531] = 8'h04 ;
            rom[5532] = 8'h1a ;
            rom[5533] = 8'h1a ;
            rom[5534] = 8'hef ;
            rom[5535] = 8'hfb ;
            rom[5536] = 8'h0d ;
            rom[5537] = 8'h04 ;
            rom[5538] = 8'hb3 ;
            rom[5539] = 8'h0b ;
            rom[5540] = 8'hd9 ;
            rom[5541] = 8'h12 ;
            rom[5542] = 8'h02 ;
            rom[5543] = 8'h16 ;
            rom[5544] = 8'hff ;
            rom[5545] = 8'he8 ;
            rom[5546] = 8'h11 ;
            rom[5547] = 8'hd9 ;
            rom[5548] = 8'he9 ;
            rom[5549] = 8'hec ;
            rom[5550] = 8'h19 ;
            rom[5551] = 8'h0e ;
            rom[5552] = 8'he8 ;
            rom[5553] = 8'hd9 ;
            rom[5554] = 8'h05 ;
            rom[5555] = 8'hee ;
            rom[5556] = 8'hf8 ;
            rom[5557] = 8'h0d ;
            rom[5558] = 8'heb ;
            rom[5559] = 8'hf3 ;
            rom[5560] = 8'hf7 ;
            rom[5561] = 8'h11 ;
            rom[5562] = 8'he7 ;
            rom[5563] = 8'hfc ;
            rom[5564] = 8'h0e ;
            rom[5565] = 8'hf8 ;
            rom[5566] = 8'h12 ;
            rom[5567] = 8'he7 ;
            rom[5568] = 8'h03 ;
            rom[5569] = 8'hc1 ;
            rom[5570] = 8'h16 ;
            rom[5571] = 8'heb ;
            rom[5572] = 8'hf3 ;
            rom[5573] = 8'hf2 ;
            rom[5574] = 8'he5 ;
            rom[5575] = 8'heb ;
            rom[5576] = 8'hfe ;
            rom[5577] = 8'hf9 ;
            rom[5578] = 8'heb ;
            rom[5579] = 8'h0b ;
            rom[5580] = 8'h01 ;
            rom[5581] = 8'h15 ;
            rom[5582] = 8'hf6 ;
            rom[5583] = 8'h1c ;
            rom[5584] = 8'h1b ;
            rom[5585] = 8'hfb ;
            rom[5586] = 8'hd4 ;
            rom[5587] = 8'h1b ;
            rom[5588] = 8'hf3 ;
            rom[5589] = 8'hf1 ;
            rom[5590] = 8'hfe ;
            rom[5591] = 8'h16 ;
            rom[5592] = 8'h15 ;
            rom[5593] = 8'h09 ;
            rom[5594] = 8'hed ;
            rom[5595] = 8'h0c ;
            rom[5596] = 8'h12 ;
            rom[5597] = 8'hd8 ;
            rom[5598] = 8'he3 ;
            rom[5599] = 8'h10 ;
            rom[5600] = 8'h07 ;
            rom[5601] = 8'h11 ;
            rom[5602] = 8'hf4 ;
            rom[5603] = 8'h0b ;
            rom[5604] = 8'hec ;
            rom[5605] = 8'hf7 ;
            rom[5606] = 8'h08 ;
            rom[5607] = 8'h0a ;
            rom[5608] = 8'hf8 ;
            rom[5609] = 8'h0c ;
            rom[5610] = 8'h1d ;
            rom[5611] = 8'hc4 ;
            rom[5612] = 8'h04 ;
            rom[5613] = 8'h0b ;
            rom[5614] = 8'h0e ;
            rom[5615] = 8'hf2 ;
            rom[5616] = 8'he5 ;
            rom[5617] = 8'h07 ;
            rom[5618] = 8'h0b ;
            rom[5619] = 8'hf5 ;
            rom[5620] = 8'h1f ;
            rom[5621] = 8'hf4 ;
            rom[5622] = 8'h07 ;
            rom[5623] = 8'h04 ;
            rom[5624] = 8'hf3 ;
            rom[5625] = 8'hed ;
            rom[5626] = 8'h0a ;
            rom[5627] = 8'hec ;
            rom[5628] = 8'h0c ;
            rom[5629] = 8'h1a ;
            rom[5630] = 8'hfa ;
            rom[5631] = 8'hf8 ;
            rom[5632] = 8'h06 ;
            rom[5633] = 8'he4 ;
            rom[5634] = 8'hdf ;
            rom[5635] = 8'hfd ;
            rom[5636] = 8'hf7 ;
            rom[5637] = 8'hfa ;
            rom[5638] = 8'hfc ;
            rom[5639] = 8'h0e ;
            rom[5640] = 8'h1d ;
            rom[5641] = 8'h08 ;
            rom[5642] = 8'hd3 ;
            rom[5643] = 8'he5 ;
            rom[5644] = 8'hf1 ;
            rom[5645] = 8'hea ;
            rom[5646] = 8'heb ;
            rom[5647] = 8'h0d ;
            rom[5648] = 8'hef ;
            rom[5649] = 8'hf8 ;
            rom[5650] = 8'h02 ;
            rom[5651] = 8'h01 ;
            rom[5652] = 8'hf8 ;
            rom[5653] = 8'he1 ;
            rom[5654] = 8'h1e ;
            rom[5655] = 8'hea ;
            rom[5656] = 8'h15 ;
            rom[5657] = 8'h1d ;
            rom[5658] = 8'h00 ;
            rom[5659] = 8'hfc ;
            rom[5660] = 8'h05 ;
            rom[5661] = 8'h06 ;
            rom[5662] = 8'h08 ;
            rom[5663] = 8'hec ;
            rom[5664] = 8'hfe ;
            rom[5665] = 8'hd5 ;
            rom[5666] = 8'h04 ;
            rom[5667] = 8'h19 ;
            rom[5668] = 8'hf6 ;
            rom[5669] = 8'hf8 ;
            rom[5670] = 8'hfc ;
            rom[5671] = 8'hf8 ;
            rom[5672] = 8'h16 ;
            rom[5673] = 8'hed ;
            rom[5674] = 8'hfc ;
            rom[5675] = 8'hff ;
            rom[5676] = 8'hfa ;
            rom[5677] = 8'hff ;
            rom[5678] = 8'hfd ;
            rom[5679] = 8'h0d ;
            rom[5680] = 8'h01 ;
            rom[5681] = 8'hfb ;
            rom[5682] = 8'hf3 ;
            rom[5683] = 8'h17 ;
            rom[5684] = 8'hea ;
            rom[5685] = 8'hf5 ;
            rom[5686] = 8'he2 ;
            rom[5687] = 8'hd7 ;
            rom[5688] = 8'h0a ;
            rom[5689] = 8'hfc ;
            rom[5690] = 8'he8 ;
            rom[5691] = 8'h0b ;
            rom[5692] = 8'h1c ;
            rom[5693] = 8'h03 ;
            rom[5694] = 8'hee ;
            rom[5695] = 8'hed ;
            rom[5696] = 8'he0 ;
            rom[5697] = 8'h05 ;
            rom[5698] = 8'he4 ;
            rom[5699] = 8'h0f ;
            rom[5700] = 8'hfa ;
            rom[5701] = 8'h01 ;
            rom[5702] = 8'h15 ;
            rom[5703] = 8'h04 ;
            rom[5704] = 8'h0d ;
            rom[5705] = 8'h03 ;
            rom[5706] = 8'ha6 ;
            rom[5707] = 8'hf2 ;
            rom[5708] = 8'hd0 ;
            rom[5709] = 8'hf2 ;
            rom[5710] = 8'h07 ;
            rom[5711] = 8'h0c ;
            rom[5712] = 8'h1c ;
            rom[5713] = 8'hfd ;
            rom[5714] = 8'hf9 ;
            rom[5715] = 8'hf2 ;
            rom[5716] = 8'h09 ;
            rom[5717] = 8'h13 ;
            rom[5718] = 8'h09 ;
            rom[5719] = 8'h01 ;
            rom[5720] = 8'hef ;
            rom[5721] = 8'h08 ;
            rom[5722] = 8'h02 ;
            rom[5723] = 8'h25 ;
            rom[5724] = 8'hfd ;
            rom[5725] = 8'hf8 ;
            rom[5726] = 8'h12 ;
            rom[5727] = 8'he4 ;
            rom[5728] = 8'hfa ;
            rom[5729] = 8'hfe ;
            rom[5730] = 8'h1a ;
            rom[5731] = 8'h08 ;
            rom[5732] = 8'he9 ;
            rom[5733] = 8'h00 ;
            rom[5734] = 8'heb ;
            rom[5735] = 8'hfc ;
            rom[5736] = 8'h20 ;
            rom[5737] = 8'hfe ;
            rom[5738] = 8'he6 ;
            rom[5739] = 8'hdb ;
            rom[5740] = 8'hea ;
            rom[5741] = 8'hf7 ;
            rom[5742] = 8'he3 ;
            rom[5743] = 8'hfe ;
            rom[5744] = 8'h02 ;
            rom[5745] = 8'h18 ;
            rom[5746] = 8'hf3 ;
            rom[5747] = 8'h09 ;
            rom[5748] = 8'h03 ;
            rom[5749] = 8'h07 ;
            rom[5750] = 8'hf5 ;
            rom[5751] = 8'h09 ;
            rom[5752] = 8'he3 ;
            rom[5753] = 8'h18 ;
            rom[5754] = 8'hf4 ;
            rom[5755] = 8'hf6 ;
            rom[5756] = 8'hfb ;
            rom[5757] = 8'h08 ;
            rom[5758] = 8'h08 ;
            rom[5759] = 8'h04 ;
            rom[5760] = 8'hfe ;
            rom[5761] = 8'h0d ;
            rom[5762] = 8'h01 ;
            rom[5763] = 8'he6 ;
            rom[5764] = 8'hf6 ;
            rom[5765] = 8'h02 ;
            rom[5766] = 8'hff ;
            rom[5767] = 8'h03 ;
            rom[5768] = 8'h08 ;
            rom[5769] = 8'hf3 ;
            rom[5770] = 8'he3 ;
            rom[5771] = 8'hfd ;
            rom[5772] = 8'h0e ;
            rom[5773] = 8'hff ;
            rom[5774] = 8'hfb ;
            rom[5775] = 8'h1f ;
            rom[5776] = 8'h0d ;
            rom[5777] = 8'h0c ;
            rom[5778] = 8'h05 ;
            rom[5779] = 8'hf0 ;
            rom[5780] = 8'he8 ;
            rom[5781] = 8'h00 ;
            rom[5782] = 8'h0f ;
            rom[5783] = 8'h14 ;
            rom[5784] = 8'hf9 ;
            rom[5785] = 8'h1b ;
            rom[5786] = 8'h10 ;
            rom[5787] = 8'h23 ;
            rom[5788] = 8'h03 ;
            rom[5789] = 8'hfb ;
            rom[5790] = 8'h03 ;
            rom[5791] = 8'hfa ;
            rom[5792] = 8'h11 ;
            rom[5793] = 8'hf7 ;
            rom[5794] = 8'h1a ;
            rom[5795] = 8'h0b ;
            rom[5796] = 8'hec ;
            rom[5797] = 8'h0e ;
            rom[5798] = 8'hef ;
            rom[5799] = 8'h00 ;
            rom[5800] = 8'h06 ;
            rom[5801] = 8'h1c ;
            rom[5802] = 8'h0a ;
            rom[5803] = 8'hc9 ;
            rom[5804] = 8'h03 ;
            rom[5805] = 8'hf2 ;
            rom[5806] = 8'hea ;
            rom[5807] = 8'hfe ;
            rom[5808] = 8'h13 ;
            rom[5809] = 8'he6 ;
            rom[5810] = 8'hdd ;
            rom[5811] = 8'h09 ;
            rom[5812] = 8'h0d ;
            rom[5813] = 8'hff ;
            rom[5814] = 8'h02 ;
            rom[5815] = 8'hfe ;
            rom[5816] = 8'hfc ;
            rom[5817] = 8'hec ;
            rom[5818] = 8'hec ;
            rom[5819] = 8'h06 ;
            rom[5820] = 8'h0d ;
            rom[5821] = 8'h1a ;
            rom[5822] = 8'h04 ;
            rom[5823] = 8'h05 ;
            rom[5824] = 8'hf0 ;
            rom[5825] = 8'hf3 ;
            rom[5826] = 8'h11 ;
            rom[5827] = 8'he1 ;
            rom[5828] = 8'hef ;
            rom[5829] = 8'heb ;
            rom[5830] = 8'he8 ;
            rom[5831] = 8'h02 ;
            rom[5832] = 8'h0d ;
            rom[5833] = 8'h15 ;
            rom[5834] = 8'hd3 ;
            rom[5835] = 8'h0d ;
            rom[5836] = 8'hf7 ;
            rom[5837] = 8'h10 ;
            rom[5838] = 8'hff ;
            rom[5839] = 8'h34 ;
            rom[5840] = 8'h1a ;
            rom[5841] = 8'h04 ;
            rom[5842] = 8'he5 ;
            rom[5843] = 8'h18 ;
            rom[5844] = 8'heb ;
            rom[5845] = 8'h06 ;
            rom[5846] = 8'hfe ;
            rom[5847] = 8'h0a ;
            rom[5848] = 8'h12 ;
            rom[5849] = 8'h06 ;
            rom[5850] = 8'hf7 ;
            rom[5851] = 8'h0e ;
            rom[5852] = 8'h18 ;
            rom[5853] = 8'he6 ;
            rom[5854] = 8'hf8 ;
            rom[5855] = 8'hfb ;
            rom[5856] = 8'h0b ;
            rom[5857] = 8'he1 ;
            rom[5858] = 8'he6 ;
            rom[5859] = 8'he4 ;
            rom[5860] = 8'hf3 ;
            rom[5861] = 8'hf8 ;
            rom[5862] = 8'h07 ;
            rom[5863] = 8'heb ;
            rom[5864] = 8'h02 ;
            rom[5865] = 8'h1b ;
            rom[5866] = 8'hfa ;
            rom[5867] = 8'hd4 ;
            rom[5868] = 8'hf9 ;
            rom[5869] = 8'hff ;
            rom[5870] = 8'hf2 ;
            rom[5871] = 8'h06 ;
            rom[5872] = 8'heb ;
            rom[5873] = 8'hf4 ;
            rom[5874] = 8'h06 ;
            rom[5875] = 8'hef ;
            rom[5876] = 8'h16 ;
            rom[5877] = 8'h00 ;
            rom[5878] = 8'hf7 ;
            rom[5879] = 8'hf9 ;
            rom[5880] = 8'h01 ;
            rom[5881] = 8'he7 ;
            rom[5882] = 8'hf0 ;
            rom[5883] = 8'hf3 ;
            rom[5884] = 8'h1d ;
            rom[5885] = 8'hfb ;
            rom[5886] = 8'h17 ;
            rom[5887] = 8'hea ;
            rom[5888] = 8'h00 ;
            rom[5889] = 8'hdd ;
            rom[5890] = 8'h20 ;
            rom[5891] = 8'h1b ;
            rom[5892] = 8'h12 ;
            rom[5893] = 8'hdb ;
            rom[5894] = 8'hd5 ;
            rom[5895] = 8'hf5 ;
            rom[5896] = 8'h0c ;
            rom[5897] = 8'h15 ;
            rom[5898] = 8'hf4 ;
            rom[5899] = 8'h0b ;
            rom[5900] = 8'hf1 ;
            rom[5901] = 8'he6 ;
            rom[5902] = 8'h01 ;
            rom[5903] = 8'hf8 ;
            rom[5904] = 8'h04 ;
            rom[5905] = 8'h32 ;
            rom[5906] = 8'he6 ;
            rom[5907] = 8'h0a ;
            rom[5908] = 8'h15 ;
            rom[5909] = 8'h17 ;
            rom[5910] = 8'h11 ;
            rom[5911] = 8'h10 ;
            rom[5912] = 8'h02 ;
            rom[5913] = 8'h25 ;
            rom[5914] = 8'hfa ;
            rom[5915] = 8'hfd ;
            rom[5916] = 8'h1e ;
            rom[5917] = 8'hf9 ;
            rom[5918] = 8'hd4 ;
            rom[5919] = 8'hef ;
            rom[5920] = 8'h13 ;
            rom[5921] = 8'hfc ;
            rom[5922] = 8'hec ;
            rom[5923] = 8'h0c ;
            rom[5924] = 8'hfe ;
            rom[5925] = 8'hf2 ;
            rom[5926] = 8'h15 ;
            rom[5927] = 8'he0 ;
            rom[5928] = 8'hf8 ;
            rom[5929] = 8'h05 ;
            rom[5930] = 8'h1d ;
            rom[5931] = 8'h06 ;
            rom[5932] = 8'h03 ;
            rom[5933] = 8'hed ;
            rom[5934] = 8'h10 ;
            rom[5935] = 8'h04 ;
            rom[5936] = 8'h1c ;
            rom[5937] = 8'hf9 ;
            rom[5938] = 8'h34 ;
            rom[5939] = 8'h02 ;
            rom[5940] = 8'h05 ;
            rom[5941] = 8'hdf ;
            rom[5942] = 8'h0a ;
            rom[5943] = 8'h0b ;
            rom[5944] = 8'hf6 ;
            rom[5945] = 8'he4 ;
            rom[5946] = 8'h06 ;
            rom[5947] = 8'he0 ;
            rom[5948] = 8'h08 ;
            rom[5949] = 8'h19 ;
            rom[5950] = 8'h10 ;
            rom[5951] = 8'hfd ;
            rom[5952] = 8'h17 ;
            rom[5953] = 8'h02 ;
            rom[5954] = 8'he1 ;
            rom[5955] = 8'hf8 ;
            rom[5956] = 8'h0b ;
            rom[5957] = 8'h0d ;
            rom[5958] = 8'h0a ;
            rom[5959] = 8'he7 ;
            rom[5960] = 8'h08 ;
            rom[5961] = 8'h0b ;
            rom[5962] = 8'h05 ;
            rom[5963] = 8'h17 ;
            rom[5964] = 8'h04 ;
            rom[5965] = 8'he9 ;
            rom[5966] = 8'h18 ;
            rom[5967] = 8'h05 ;
            rom[5968] = 8'h0f ;
            rom[5969] = 8'hef ;
            rom[5970] = 8'h1f ;
            rom[5971] = 8'h0f ;
            rom[5972] = 8'h1c ;
            rom[5973] = 8'hff ;
            rom[5974] = 8'hfa ;
            rom[5975] = 8'hee ;
            rom[5976] = 8'h09 ;
            rom[5977] = 8'h13 ;
            rom[5978] = 8'hfb ;
            rom[5979] = 8'h26 ;
            rom[5980] = 8'h0a ;
            rom[5981] = 8'h03 ;
            rom[5982] = 8'hf3 ;
            rom[5983] = 8'h0a ;
            rom[5984] = 8'h1a ;
            rom[5985] = 8'hf7 ;
            rom[5986] = 8'h0d ;
            rom[5987] = 8'h29 ;
            rom[5988] = 8'h1a ;
            rom[5989] = 8'h08 ;
            rom[5990] = 8'hf2 ;
            rom[5991] = 8'hcd ;
            rom[5992] = 8'heb ;
            rom[5993] = 8'hdf ;
            rom[5994] = 8'hf0 ;
            rom[5995] = 8'hed ;
            rom[5996] = 8'h08 ;
            rom[5997] = 8'hed ;
            rom[5998] = 8'h09 ;
            rom[5999] = 8'he4 ;
            rom[6000] = 8'h0b ;
            rom[6001] = 8'hef ;
            rom[6002] = 8'h11 ;
            rom[6003] = 8'h22 ;
            rom[6004] = 8'hef ;
            rom[6005] = 8'h05 ;
            rom[6006] = 8'hf7 ;
            rom[6007] = 8'hea ;
            rom[6008] = 8'hfa ;
            rom[6009] = 8'hf4 ;
            rom[6010] = 8'h06 ;
            rom[6011] = 8'h0e ;
            rom[6012] = 8'h1f ;
            rom[6013] = 8'he3 ;
            rom[6014] = 8'hd7 ;
            rom[6015] = 8'he7 ;
            rom[6016] = 8'he5 ;
            rom[6017] = 8'h02 ;
            rom[6018] = 8'h01 ;
            rom[6019] = 8'h10 ;
            rom[6020] = 8'he7 ;
            rom[6021] = 8'h01 ;
            rom[6022] = 8'h0b ;
            rom[6023] = 8'he9 ;
            rom[6024] = 8'h11 ;
            rom[6025] = 8'h22 ;
            rom[6026] = 8'h01 ;
            rom[6027] = 8'hfc ;
            rom[6028] = 8'h0f ;
            rom[6029] = 8'hee ;
            rom[6030] = 8'h0c ;
            rom[6031] = 8'h01 ;
            rom[6032] = 8'hef ;
            rom[6033] = 8'hf7 ;
            rom[6034] = 8'hfb ;
            rom[6035] = 8'hfa ;
            rom[6036] = 8'h27 ;
            rom[6037] = 8'hc5 ;
            rom[6038] = 8'h1a ;
            rom[6039] = 8'h00 ;
            rom[6040] = 8'hbc ;
            rom[6041] = 8'hfe ;
            rom[6042] = 8'hff ;
            rom[6043] = 8'h0b ;
            rom[6044] = 8'hf9 ;
            rom[6045] = 8'h10 ;
            rom[6046] = 8'h01 ;
            rom[6047] = 8'h0d ;
            rom[6048] = 8'h03 ;
            rom[6049] = 8'h04 ;
            rom[6050] = 8'h02 ;
            rom[6051] = 8'hf0 ;
            rom[6052] = 8'hf8 ;
            rom[6053] = 8'hfb ;
            rom[6054] = 8'hf8 ;
            rom[6055] = 8'h2a ;
            rom[6056] = 8'hf9 ;
            rom[6057] = 8'hf0 ;
            rom[6058] = 8'h11 ;
            rom[6059] = 8'h10 ;
            rom[6060] = 8'hef ;
            rom[6061] = 8'hd2 ;
            rom[6062] = 8'hee ;
            rom[6063] = 8'hf1 ;
            rom[6064] = 8'h2c ;
            rom[6065] = 8'hfc ;
            rom[6066] = 8'h00 ;
            rom[6067] = 8'hf0 ;
            rom[6068] = 8'hf2 ;
            rom[6069] = 8'hd6 ;
            rom[6070] = 8'h00 ;
            rom[6071] = 8'hf5 ;
            rom[6072] = 8'h09 ;
            rom[6073] = 8'h14 ;
            rom[6074] = 8'he2 ;
            rom[6075] = 8'h09 ;
            rom[6076] = 8'hfe ;
            rom[6077] = 8'hf6 ;
            rom[6078] = 8'hf4 ;
            rom[6079] = 8'he9 ;
            rom[6080] = 8'h1b ;
            rom[6081] = 8'hf9 ;
            rom[6082] = 8'h0c ;
            rom[6083] = 8'h17 ;
            rom[6084] = 8'hf6 ;
            rom[6085] = 8'h0c ;
            rom[6086] = 8'h05 ;
            rom[6087] = 8'h00 ;
            rom[6088] = 8'h12 ;
            rom[6089] = 8'h06 ;
            rom[6090] = 8'h1f ;
            rom[6091] = 8'h09 ;
            rom[6092] = 8'h23 ;
            rom[6093] = 8'h07 ;
            rom[6094] = 8'h09 ;
            rom[6095] = 8'he9 ;
            rom[6096] = 8'h08 ;
            rom[6097] = 8'he2 ;
            rom[6098] = 8'hea ;
            rom[6099] = 8'h1c ;
            rom[6100] = 8'hf0 ;
            rom[6101] = 8'hec ;
            rom[6102] = 8'h06 ;
            rom[6103] = 8'hfe ;
            rom[6104] = 8'h22 ;
            rom[6105] = 8'h02 ;
            rom[6106] = 8'hfd ;
            rom[6107] = 8'h17 ;
            rom[6108] = 8'hfd ;
            rom[6109] = 8'hef ;
            rom[6110] = 8'hef ;
            rom[6111] = 8'h1a ;
            rom[6112] = 8'hfa ;
            rom[6113] = 8'h0c ;
            rom[6114] = 8'h2d ;
            rom[6115] = 8'h14 ;
            rom[6116] = 8'h07 ;
            rom[6117] = 8'h18 ;
            rom[6118] = 8'hee ;
            rom[6119] = 8'hb4 ;
            rom[6120] = 8'he3 ;
            rom[6121] = 8'h11 ;
            rom[6122] = 8'hf6 ;
            rom[6123] = 8'hf1 ;
            rom[6124] = 8'h11 ;
            rom[6125] = 8'h05 ;
            rom[6126] = 8'he9 ;
            rom[6127] = 8'h03 ;
            rom[6128] = 8'hf0 ;
            rom[6129] = 8'h0a ;
            rom[6130] = 8'hf8 ;
            rom[6131] = 8'h15 ;
            rom[6132] = 8'hf2 ;
            rom[6133] = 8'hed ;
            rom[6134] = 8'h0e ;
            rom[6135] = 8'h0d ;
            rom[6136] = 8'hf6 ;
            rom[6137] = 8'h03 ;
            rom[6138] = 8'hdd ;
            rom[6139] = 8'h18 ;
            rom[6140] = 8'hf5 ;
            rom[6141] = 8'hef ;
            rom[6142] = 8'hff ;
            rom[6143] = 8'h13 ;
            rom[6144] = 8'h18 ;
            rom[6145] = 8'hff ;
            rom[6146] = 8'hf2 ;
            rom[6147] = 8'hf4 ;
            rom[6148] = 8'hfe ;
            rom[6149] = 8'hfb ;
            rom[6150] = 8'hf4 ;
            rom[6151] = 8'hb3 ;
            rom[6152] = 8'hf5 ;
            rom[6153] = 8'hfa ;
            rom[6154] = 8'h06 ;
            rom[6155] = 8'h06 ;
            rom[6156] = 8'hd4 ;
            rom[6157] = 8'he1 ;
            rom[6158] = 8'h03 ;
            rom[6159] = 8'hef ;
            rom[6160] = 8'heb ;
            rom[6161] = 8'he6 ;
            rom[6162] = 8'hf8 ;
            rom[6163] = 8'hf6 ;
            rom[6164] = 8'hda ;
            rom[6165] = 8'h15 ;
            rom[6166] = 8'h09 ;
            rom[6167] = 8'h03 ;
            rom[6168] = 8'hee ;
            rom[6169] = 8'hf7 ;
            rom[6170] = 8'h0d ;
            rom[6171] = 8'hd8 ;
            rom[6172] = 8'hfc ;
            rom[6173] = 8'hed ;
            rom[6174] = 8'hde ;
            rom[6175] = 8'hf7 ;
            rom[6176] = 8'h08 ;
            rom[6177] = 8'h03 ;
            rom[6178] = 8'hfd ;
            rom[6179] = 8'h00 ;
            rom[6180] = 8'hd7 ;
            rom[6181] = 8'hfc ;
            rom[6182] = 8'hf2 ;
            rom[6183] = 8'h07 ;
            rom[6184] = 8'hef ;
            rom[6185] = 8'hff ;
            rom[6186] = 8'he3 ;
            rom[6187] = 8'hfa ;
            rom[6188] = 8'h05 ;
            rom[6189] = 8'hf3 ;
            rom[6190] = 8'h00 ;
            rom[6191] = 8'hd5 ;
            rom[6192] = 8'hef ;
            rom[6193] = 8'h16 ;
            rom[6194] = 8'hf7 ;
            rom[6195] = 8'he3 ;
            rom[6196] = 8'hf0 ;
            rom[6197] = 8'h09 ;
            rom[6198] = 8'hf1 ;
            rom[6199] = 8'h0c ;
            rom[6200] = 8'h11 ;
            rom[6201] = 8'h0e ;
            rom[6202] = 8'hdf ;
            rom[6203] = 8'hde ;
            rom[6204] = 8'hff ;
            rom[6205] = 8'h12 ;
            rom[6206] = 8'h02 ;
            rom[6207] = 8'hf5 ;
            rom[6208] = 8'h0f ;
            rom[6209] = 8'he8 ;
            rom[6210] = 8'h12 ;
            rom[6211] = 8'h06 ;
            rom[6212] = 8'h1e ;
            rom[6213] = 8'hf4 ;
            rom[6214] = 8'hf4 ;
            rom[6215] = 8'heb ;
            rom[6216] = 8'hdb ;
            rom[6217] = 8'hfe ;
            rom[6218] = 8'hfb ;
            rom[6219] = 8'hfa ;
            rom[6220] = 8'hf4 ;
            rom[6221] = 8'hff ;
            rom[6222] = 8'hf7 ;
            rom[6223] = 8'hf7 ;
            rom[6224] = 8'hfa ;
            rom[6225] = 8'h0c ;
            rom[6226] = 8'h03 ;
            rom[6227] = 8'h23 ;
            rom[6228] = 8'he8 ;
            rom[6229] = 8'hf7 ;
            rom[6230] = 8'hfe ;
            rom[6231] = 8'h01 ;
            rom[6232] = 8'h17 ;
            rom[6233] = 8'hd6 ;
            rom[6234] = 8'hff ;
            rom[6235] = 8'hee ;
            rom[6236] = 8'he8 ;
            rom[6237] = 8'hed ;
            rom[6238] = 8'h02 ;
            rom[6239] = 8'hfd ;
            rom[6240] = 8'he8 ;
            rom[6241] = 8'hf1 ;
            rom[6242] = 8'he8 ;
            rom[6243] = 8'hff ;
            rom[6244] = 8'h22 ;
            rom[6245] = 8'hf2 ;
            rom[6246] = 8'h1c ;
            rom[6247] = 8'hd2 ;
            rom[6248] = 8'h0d ;
            rom[6249] = 8'he7 ;
            rom[6250] = 8'h0f ;
            rom[6251] = 8'hfd ;
            rom[6252] = 8'h02 ;
            rom[6253] = 8'h11 ;
            rom[6254] = 8'hf6 ;
            rom[6255] = 8'h17 ;
            rom[6256] = 8'h06 ;
            rom[6257] = 8'hf1 ;
            rom[6258] = 8'h12 ;
            rom[6259] = 8'hfd ;
            rom[6260] = 8'he8 ;
            rom[6261] = 8'hf3 ;
            rom[6262] = 8'hff ;
            rom[6263] = 8'h0a ;
            rom[6264] = 8'hf8 ;
            rom[6265] = 8'he9 ;
            rom[6266] = 8'hf5 ;
            rom[6267] = 8'h0b ;
            rom[6268] = 8'h13 ;
            rom[6269] = 8'hea ;
            rom[6270] = 8'h09 ;
            rom[6271] = 8'h00 ;
            rom[6272] = 8'h07 ;
            rom[6273] = 8'hfc ;
            rom[6274] = 8'hd5 ;
            rom[6275] = 8'h09 ;
            rom[6276] = 8'h13 ;
            rom[6277] = 8'hd6 ;
            rom[6278] = 8'h0a ;
            rom[6279] = 8'h0f ;
            rom[6280] = 8'hd5 ;
            rom[6281] = 8'hd3 ;
            rom[6282] = 8'hfb ;
            rom[6283] = 8'hf7 ;
            rom[6284] = 8'hf5 ;
            rom[6285] = 8'he6 ;
            rom[6286] = 8'h10 ;
            rom[6287] = 8'hf8 ;
            rom[6288] = 8'hfb ;
            rom[6289] = 8'h09 ;
            rom[6290] = 8'hfa ;
            rom[6291] = 8'hdd ;
            rom[6292] = 8'hfb ;
            rom[6293] = 8'h14 ;
            rom[6294] = 8'h13 ;
            rom[6295] = 8'he2 ;
            rom[6296] = 8'hcf ;
            rom[6297] = 8'h05 ;
            rom[6298] = 8'he2 ;
            rom[6299] = 8'h13 ;
            rom[6300] = 8'he8 ;
            rom[6301] = 8'he0 ;
            rom[6302] = 8'hfb ;
            rom[6303] = 8'h0c ;
            rom[6304] = 8'hdc ;
            rom[6305] = 8'hed ;
            rom[6306] = 8'h03 ;
            rom[6307] = 8'h15 ;
            rom[6308] = 8'heb ;
            rom[6309] = 8'h08 ;
            rom[6310] = 8'hed ;
            rom[6311] = 8'hfd ;
            rom[6312] = 8'hdd ;
            rom[6313] = 8'h05 ;
            rom[6314] = 8'h02 ;
            rom[6315] = 8'h0c ;
            rom[6316] = 8'hff ;
            rom[6317] = 8'h09 ;
            rom[6318] = 8'h08 ;
            rom[6319] = 8'h0f ;
            rom[6320] = 8'h0b ;
            rom[6321] = 8'h0e ;
            rom[6322] = 8'hfb ;
            rom[6323] = 8'hed ;
            rom[6324] = 8'h09 ;
            rom[6325] = 8'h0a ;
            rom[6326] = 8'hf8 ;
            rom[6327] = 8'hfc ;
            rom[6328] = 8'hd1 ;
            rom[6329] = 8'hfb ;
            rom[6330] = 8'h1b ;
            rom[6331] = 8'hff ;
            rom[6332] = 8'he2 ;
            rom[6333] = 8'he8 ;
            rom[6334] = 8'h1d ;
            rom[6335] = 8'h0e ;
            rom[6336] = 8'hfe ;
            rom[6337] = 8'h15 ;
            rom[6338] = 8'hf8 ;
            rom[6339] = 8'hf7 ;
            rom[6340] = 8'h13 ;
            rom[6341] = 8'h06 ;
            rom[6342] = 8'hdb ;
            rom[6343] = 8'h00 ;
            rom[6344] = 8'he6 ;
            rom[6345] = 8'he6 ;
            rom[6346] = 8'hfb ;
            rom[6347] = 8'h1b ;
            rom[6348] = 8'he9 ;
            rom[6349] = 8'h18 ;
            rom[6350] = 8'h30 ;
            rom[6351] = 8'h10 ;
            rom[6352] = 8'hfa ;
            rom[6353] = 8'hfa ;
            rom[6354] = 8'h1d ;
            rom[6355] = 8'hf3 ;
            rom[6356] = 8'hfa ;
            rom[6357] = 8'he6 ;
            rom[6358] = 8'hfb ;
            rom[6359] = 8'he7 ;
            rom[6360] = 8'h06 ;
            rom[6361] = 8'h14 ;
            rom[6362] = 8'hf2 ;
            rom[6363] = 8'h0a ;
            rom[6364] = 8'h0a ;
            rom[6365] = 8'hf4 ;
            rom[6366] = 8'h1a ;
            rom[6367] = 8'h2e ;
            rom[6368] = 8'he8 ;
            rom[6369] = 8'hf7 ;
            rom[6370] = 8'h17 ;
            rom[6371] = 8'h0c ;
            rom[6372] = 8'h0e ;
            rom[6373] = 8'h03 ;
            rom[6374] = 8'h05 ;
            rom[6375] = 8'h0c ;
            rom[6376] = 8'he1 ;
            rom[6377] = 8'h01 ;
            rom[6378] = 8'hf5 ;
            rom[6379] = 8'h0e ;
            rom[6380] = 8'h1f ;
            rom[6381] = 8'hf2 ;
            rom[6382] = 8'hf1 ;
            rom[6383] = 8'hd0 ;
            rom[6384] = 8'h16 ;
            rom[6385] = 8'h07 ;
            rom[6386] = 8'hed ;
            rom[6387] = 8'he8 ;
            rom[6388] = 8'hf2 ;
            rom[6389] = 8'hf8 ;
            rom[6390] = 8'hee ;
            rom[6391] = 8'h14 ;
            rom[6392] = 8'hf1 ;
            rom[6393] = 8'h08 ;
            rom[6394] = 8'h1f ;
            rom[6395] = 8'he2 ;
            rom[6396] = 8'hda ;
            rom[6397] = 8'h08 ;
            rom[6398] = 8'hee ;
            rom[6399] = 8'hfd ;
            rom[6400] = 8'h21 ;
            rom[6401] = 8'hed ;
            rom[6402] = 8'h19 ;
            rom[6403] = 8'h07 ;
            rom[6404] = 8'h10 ;
            rom[6405] = 8'h11 ;
            rom[6406] = 8'h05 ;
            rom[6407] = 8'h0c ;
            rom[6408] = 8'hd9 ;
            rom[6409] = 8'hf1 ;
            rom[6410] = 8'hfd ;
            rom[6411] = 8'h05 ;
            rom[6412] = 8'he3 ;
            rom[6413] = 8'he8 ;
            rom[6414] = 8'hfe ;
            rom[6415] = 8'hf6 ;
            rom[6416] = 8'hea ;
            rom[6417] = 8'hf4 ;
            rom[6418] = 8'h00 ;
            rom[6419] = 8'h0b ;
            rom[6420] = 8'hf7 ;
            rom[6421] = 8'hef ;
            rom[6422] = 8'hf4 ;
            rom[6423] = 8'h13 ;
            rom[6424] = 8'h08 ;
            rom[6425] = 8'heb ;
            rom[6426] = 8'hd9 ;
            rom[6427] = 8'h19 ;
            rom[6428] = 8'h06 ;
            rom[6429] = 8'h07 ;
            rom[6430] = 8'h0d ;
            rom[6431] = 8'he4 ;
            rom[6432] = 8'h10 ;
            rom[6433] = 8'hfb ;
            rom[6434] = 8'he1 ;
            rom[6435] = 8'he4 ;
            rom[6436] = 8'h21 ;
            rom[6437] = 8'h2d ;
            rom[6438] = 8'hec ;
            rom[6439] = 8'he5 ;
            rom[6440] = 8'h14 ;
            rom[6441] = 8'hb1 ;
            rom[6442] = 8'he5 ;
            rom[6443] = 8'hff ;
            rom[6444] = 8'hd6 ;
            rom[6445] = 8'h18 ;
            rom[6446] = 8'hc4 ;
            rom[6447] = 8'h1c ;
            rom[6448] = 8'hf8 ;
            rom[6449] = 8'h16 ;
            rom[6450] = 8'h1f ;
            rom[6451] = 8'hf7 ;
            rom[6452] = 8'hf8 ;
            rom[6453] = 8'hf9 ;
            rom[6454] = 8'hea ;
            rom[6455] = 8'h03 ;
            rom[6456] = 8'h04 ;
            rom[6457] = 8'hf2 ;
            rom[6458] = 8'heb ;
            rom[6459] = 8'h06 ;
            rom[6460] = 8'hf4 ;
            rom[6461] = 8'hf9 ;
            rom[6462] = 8'he8 ;
            rom[6463] = 8'h02 ;
            rom[6464] = 8'h16 ;
            rom[6465] = 8'h12 ;
            rom[6466] = 8'hf9 ;
            rom[6467] = 8'h02 ;
            rom[6468] = 8'h19 ;
            rom[6469] = 8'hef ;
            rom[6470] = 8'h04 ;
            rom[6471] = 8'h10 ;
            rom[6472] = 8'h18 ;
            rom[6473] = 8'hc9 ;
            rom[6474] = 8'h0f ;
            rom[6475] = 8'h07 ;
            rom[6476] = 8'h19 ;
            rom[6477] = 8'h07 ;
            rom[6478] = 8'hf6 ;
            rom[6479] = 8'hfc ;
            rom[6480] = 8'h16 ;
            rom[6481] = 8'h0c ;
            rom[6482] = 8'hdf ;
            rom[6483] = 8'he3 ;
            rom[6484] = 8'hf9 ;
            rom[6485] = 8'hf6 ;
            rom[6486] = 8'hdb ;
            rom[6487] = 8'h19 ;
            rom[6488] = 8'hf7 ;
            rom[6489] = 8'hd3 ;
            rom[6490] = 8'hed ;
            rom[6491] = 8'hf8 ;
            rom[6492] = 8'hff ;
            rom[6493] = 8'h08 ;
            rom[6494] = 8'h18 ;
            rom[6495] = 8'h0d ;
            rom[6496] = 8'h03 ;
            rom[6497] = 8'h12 ;
            rom[6498] = 8'he7 ;
            rom[6499] = 8'hef ;
            rom[6500] = 8'h06 ;
            rom[6501] = 8'h0a ;
            rom[6502] = 8'hec ;
            rom[6503] = 8'h28 ;
            rom[6504] = 8'he7 ;
            rom[6505] = 8'hf9 ;
            rom[6506] = 8'h03 ;
            rom[6507] = 8'hf6 ;
            rom[6508] = 8'hfb ;
            rom[6509] = 8'hdc ;
            rom[6510] = 8'h14 ;
            rom[6511] = 8'he4 ;
            rom[6512] = 8'h09 ;
            rom[6513] = 8'hf9 ;
            rom[6514] = 8'hec ;
            rom[6515] = 8'h08 ;
            rom[6516] = 8'hce ;
            rom[6517] = 8'hff ;
            rom[6518] = 8'h0e ;
            rom[6519] = 8'h1f ;
            rom[6520] = 8'h03 ;
            rom[6521] = 8'hf5 ;
            rom[6522] = 8'h0d ;
            rom[6523] = 8'h10 ;
            rom[6524] = 8'hfc ;
            rom[6525] = 8'hcb ;
            rom[6526] = 8'h13 ;
            rom[6527] = 8'hf4 ;
            rom[6528] = 8'h03 ;
            rom[6529] = 8'hf6 ;
            rom[6530] = 8'hec ;
            rom[6531] = 8'hf5 ;
            rom[6532] = 8'h13 ;
            rom[6533] = 8'h0b ;
            rom[6534] = 8'h07 ;
            rom[6535] = 8'hf4 ;
            rom[6536] = 8'hd7 ;
            rom[6537] = 8'hed ;
            rom[6538] = 8'h02 ;
            rom[6539] = 8'hf9 ;
            rom[6540] = 8'hf4 ;
            rom[6541] = 8'h23 ;
            rom[6542] = 8'hf6 ;
            rom[6543] = 8'h01 ;
            rom[6544] = 8'h02 ;
            rom[6545] = 8'h1b ;
            rom[6546] = 8'h14 ;
            rom[6547] = 8'h0c ;
            rom[6548] = 8'h10 ;
            rom[6549] = 8'h0a ;
            rom[6550] = 8'h04 ;
            rom[6551] = 8'hf1 ;
            rom[6552] = 8'he1 ;
            rom[6553] = 8'hed ;
            rom[6554] = 8'h1a ;
            rom[6555] = 8'h1d ;
            rom[6556] = 8'hbf ;
            rom[6557] = 8'hfc ;
            rom[6558] = 8'hfe ;
            rom[6559] = 8'h10 ;
            rom[6560] = 8'hd9 ;
            rom[6561] = 8'hec ;
            rom[6562] = 8'h0d ;
            rom[6563] = 8'hf9 ;
            rom[6564] = 8'h11 ;
            rom[6565] = 8'h34 ;
            rom[6566] = 8'hed ;
            rom[6567] = 8'h10 ;
            rom[6568] = 8'hfc ;
            rom[6569] = 8'hff ;
            rom[6570] = 8'h08 ;
            rom[6571] = 8'h09 ;
            rom[6572] = 8'h17 ;
            rom[6573] = 8'hf5 ;
            rom[6574] = 8'hed ;
            rom[6575] = 8'hfe ;
            rom[6576] = 8'h09 ;
            rom[6577] = 8'h14 ;
            rom[6578] = 8'hd9 ;
            rom[6579] = 8'h23 ;
            rom[6580] = 8'hfa ;
            rom[6581] = 8'he9 ;
            rom[6582] = 8'hf8 ;
            rom[6583] = 8'h13 ;
            rom[6584] = 8'hdb ;
            rom[6585] = 8'hf9 ;
            rom[6586] = 8'hfb ;
            rom[6587] = 8'h25 ;
            rom[6588] = 8'hbd ;
            rom[6589] = 8'he4 ;
            rom[6590] = 8'h15 ;
            rom[6591] = 8'h1e ;
            rom[6592] = 8'hfa ;
            rom[6593] = 8'hf3 ;
            rom[6594] = 8'hfb ;
            rom[6595] = 8'heb ;
            rom[6596] = 8'h01 ;
            rom[6597] = 8'h32 ;
            rom[6598] = 8'hd7 ;
            rom[6599] = 8'hdb ;
            rom[6600] = 8'he3 ;
            rom[6601] = 8'hf5 ;
            rom[6602] = 8'h0f ;
            rom[6603] = 8'he8 ;
            rom[6604] = 8'h09 ;
            rom[6605] = 8'hee ;
            rom[6606] = 8'hf6 ;
            rom[6607] = 8'h0a ;
            rom[6608] = 8'hf5 ;
            rom[6609] = 8'h18 ;
            rom[6610] = 8'h0b ;
            rom[6611] = 8'hf1 ;
            rom[6612] = 8'h09 ;
            rom[6613] = 8'h10 ;
            rom[6614] = 8'hfa ;
            rom[6615] = 8'h21 ;
            rom[6616] = 8'hf1 ;
            rom[6617] = 8'hf8 ;
            rom[6618] = 8'hff ;
            rom[6619] = 8'hec ;
            rom[6620] = 8'h17 ;
            rom[6621] = 8'hee ;
            rom[6622] = 8'hff ;
            rom[6623] = 8'h0e ;
            rom[6624] = 8'h17 ;
            rom[6625] = 8'hf0 ;
            rom[6626] = 8'hfa ;
            rom[6627] = 8'h02 ;
            rom[6628] = 8'h14 ;
            rom[6629] = 8'h2d ;
            rom[6630] = 8'h32 ;
            rom[6631] = 8'h0b ;
            rom[6632] = 8'h10 ;
            rom[6633] = 8'hf5 ;
            rom[6634] = 8'hfa ;
            rom[6635] = 8'h10 ;
            rom[6636] = 8'h2c ;
            rom[6637] = 8'h0a ;
            rom[6638] = 8'hfa ;
            rom[6639] = 8'he9 ;
            rom[6640] = 8'hfc ;
            rom[6641] = 8'hf3 ;
            rom[6642] = 8'h0e ;
            rom[6643] = 8'hf3 ;
            rom[6644] = 8'h22 ;
            rom[6645] = 8'hfa ;
            rom[6646] = 8'hfe ;
            rom[6647] = 8'hff ;
            rom[6648] = 8'h0c ;
            rom[6649] = 8'h04 ;
            rom[6650] = 8'h01 ;
            rom[6651] = 8'he8 ;
            rom[6652] = 8'he5 ;
            rom[6653] = 8'hc2 ;
            rom[6654] = 8'h07 ;
            rom[6655] = 8'h06 ;
            rom[6656] = 8'h15 ;
            rom[6657] = 8'h0d ;
            rom[6658] = 8'h0d ;
            rom[6659] = 8'h0d ;
            rom[6660] = 8'h0f ;
            rom[6661] = 8'h01 ;
            rom[6662] = 8'h11 ;
            rom[6663] = 8'hfc ;
            rom[6664] = 8'hf8 ;
            rom[6665] = 8'he0 ;
            rom[6666] = 8'hf5 ;
            rom[6667] = 8'hef ;
            rom[6668] = 8'hfc ;
            rom[6669] = 8'hfc ;
            rom[6670] = 8'h01 ;
            rom[6671] = 8'hf8 ;
            rom[6672] = 8'h09 ;
            rom[6673] = 8'h00 ;
            rom[6674] = 8'h11 ;
            rom[6675] = 8'hf7 ;
            rom[6676] = 8'he2 ;
            rom[6677] = 8'h15 ;
            rom[6678] = 8'hfc ;
            rom[6679] = 8'h09 ;
            rom[6680] = 8'h27 ;
            rom[6681] = 8'hd0 ;
            rom[6682] = 8'h03 ;
            rom[6683] = 8'hef ;
            rom[6684] = 8'h02 ;
            rom[6685] = 8'hf9 ;
            rom[6686] = 8'hf1 ;
            rom[6687] = 8'hce ;
            rom[6688] = 8'h15 ;
            rom[6689] = 8'hf7 ;
            rom[6690] = 8'hee ;
            rom[6691] = 8'hfd ;
            rom[6692] = 8'h26 ;
            rom[6693] = 8'hf2 ;
            rom[6694] = 8'h01 ;
            rom[6695] = 8'h05 ;
            rom[6696] = 8'hde ;
            rom[6697] = 8'hc9 ;
            rom[6698] = 8'hfd ;
            rom[6699] = 8'hf5 ;
            rom[6700] = 8'h0a ;
            rom[6701] = 8'hf3 ;
            rom[6702] = 8'he1 ;
            rom[6703] = 8'h0b ;
            rom[6704] = 8'h05 ;
            rom[6705] = 8'hdc ;
            rom[6706] = 8'h0b ;
            rom[6707] = 8'h02 ;
            rom[6708] = 8'hf2 ;
            rom[6709] = 8'h0d ;
            rom[6710] = 8'hff ;
            rom[6711] = 8'h11 ;
            rom[6712] = 8'hdb ;
            rom[6713] = 8'h10 ;
            rom[6714] = 8'h04 ;
            rom[6715] = 8'hfa ;
            rom[6716] = 8'hfe ;
            rom[6717] = 8'hea ;
            rom[6718] = 8'h04 ;
            rom[6719] = 8'h16 ;
            rom[6720] = 8'h16 ;
            rom[6721] = 8'hff ;
            rom[6722] = 8'h0f ;
            rom[6723] = 8'h07 ;
            rom[6724] = 8'h1f ;
            rom[6725] = 8'h20 ;
            rom[6726] = 8'h16 ;
            rom[6727] = 8'h05 ;
            rom[6728] = 8'hd3 ;
            rom[6729] = 8'he9 ;
            rom[6730] = 8'h24 ;
            rom[6731] = 8'hf3 ;
            rom[6732] = 8'hfa ;
            rom[6733] = 8'h09 ;
            rom[6734] = 8'hf0 ;
            rom[6735] = 8'hc0 ;
            rom[6736] = 8'hf6 ;
            rom[6737] = 8'h0b ;
            rom[6738] = 8'hfa ;
            rom[6739] = 8'h0a ;
            rom[6740] = 8'hf6 ;
            rom[6741] = 8'hed ;
            rom[6742] = 8'hfe ;
            rom[6743] = 8'h27 ;
            rom[6744] = 8'hfe ;
            rom[6745] = 8'hc5 ;
            rom[6746] = 8'hf3 ;
            rom[6747] = 8'hca ;
            rom[6748] = 8'h08 ;
            rom[6749] = 8'h1f ;
            rom[6750] = 8'hfe ;
            rom[6751] = 8'hc6 ;
            rom[6752] = 8'hed ;
            rom[6753] = 8'hf9 ;
            rom[6754] = 8'h07 ;
            rom[6755] = 8'heb ;
            rom[6756] = 8'h1e ;
            rom[6757] = 8'h0b ;
            rom[6758] = 8'h0c ;
            rom[6759] = 8'he8 ;
            rom[6760] = 8'h1d ;
            rom[6761] = 8'hf2 ;
            rom[6762] = 8'hf7 ;
            rom[6763] = 8'h16 ;
            rom[6764] = 8'h04 ;
            rom[6765] = 8'hfe ;
            rom[6766] = 8'he3 ;
            rom[6767] = 8'h1c ;
            rom[6768] = 8'hf2 ;
            rom[6769] = 8'hd4 ;
            rom[6770] = 8'h18 ;
            rom[6771] = 8'hf2 ;
            rom[6772] = 8'he8 ;
            rom[6773] = 8'hec ;
            rom[6774] = 8'h02 ;
            rom[6775] = 8'h0b ;
            rom[6776] = 8'h0a ;
            rom[6777] = 8'hfc ;
            rom[6778] = 8'hf2 ;
            rom[6779] = 8'h0a ;
            rom[6780] = 8'h02 ;
            rom[6781] = 8'hfa ;
            rom[6782] = 8'h18 ;
            rom[6783] = 8'hf4 ;
            rom[6784] = 8'heb ;
            rom[6785] = 8'hf3 ;
            rom[6786] = 8'h03 ;
            rom[6787] = 8'h2a ;
            rom[6788] = 8'hfc ;
            rom[6789] = 8'h09 ;
            rom[6790] = 8'h06 ;
            rom[6791] = 8'hd6 ;
            rom[6792] = 8'h05 ;
            rom[6793] = 8'hed ;
            rom[6794] = 8'h14 ;
            rom[6795] = 8'h09 ;
            rom[6796] = 8'h13 ;
            rom[6797] = 8'h0b ;
            rom[6798] = 8'h07 ;
            rom[6799] = 8'he0 ;
            rom[6800] = 8'he8 ;
            rom[6801] = 8'h0f ;
            rom[6802] = 8'he3 ;
            rom[6803] = 8'h10 ;
            rom[6804] = 8'h0d ;
            rom[6805] = 8'hfe ;
            rom[6806] = 8'he2 ;
            rom[6807] = 8'hf6 ;
            rom[6808] = 8'h06 ;
            rom[6809] = 8'hff ;
            rom[6810] = 8'h05 ;
            rom[6811] = 8'hc7 ;
            rom[6812] = 8'hf4 ;
            rom[6813] = 8'h37 ;
            rom[6814] = 8'h3d ;
            rom[6815] = 8'h0c ;
            rom[6816] = 8'h08 ;
            rom[6817] = 8'hfb ;
            rom[6818] = 8'hfe ;
            rom[6819] = 8'h04 ;
            rom[6820] = 8'hf0 ;
            rom[6821] = 8'h0f ;
            rom[6822] = 8'h00 ;
            rom[6823] = 8'hf3 ;
            rom[6824] = 8'hfa ;
            rom[6825] = 8'h00 ;
            rom[6826] = 8'hda ;
            rom[6827] = 8'hff ;
            rom[6828] = 8'h47 ;
            rom[6829] = 8'hec ;
            rom[6830] = 8'h04 ;
            rom[6831] = 8'h26 ;
            rom[6832] = 8'hcf ;
            rom[6833] = 8'h02 ;
            rom[6834] = 8'h1d ;
            rom[6835] = 8'h01 ;
            rom[6836] = 8'he9 ;
            rom[6837] = 8'h11 ;
            rom[6838] = 8'h30 ;
            rom[6839] = 8'heb ;
            rom[6840] = 8'hf4 ;
            rom[6841] = 8'h02 ;
            rom[6842] = 8'h0d ;
            rom[6843] = 8'h2b ;
            rom[6844] = 8'h11 ;
            rom[6845] = 8'hef ;
            rom[6846] = 8'h16 ;
            rom[6847] = 8'h01 ;
            rom[6848] = 8'h20 ;
            rom[6849] = 8'h08 ;
            rom[6850] = 8'h07 ;
            rom[6851] = 8'h0c ;
            rom[6852] = 8'h29 ;
            rom[6853] = 8'hef ;
            rom[6854] = 8'h0a ;
            rom[6855] = 8'hfd ;
            rom[6856] = 8'hf2 ;
            rom[6857] = 8'hec ;
            rom[6858] = 8'h0a ;
            rom[6859] = 8'hfa ;
            rom[6860] = 8'h00 ;
            rom[6861] = 8'hfb ;
            rom[6862] = 8'h0a ;
            rom[6863] = 8'he4 ;
            rom[6864] = 8'h0f ;
            rom[6865] = 8'hff ;
            rom[6866] = 8'h0e ;
            rom[6867] = 8'he4 ;
            rom[6868] = 8'h0b ;
            rom[6869] = 8'h00 ;
            rom[6870] = 8'hfb ;
            rom[6871] = 8'h06 ;
            rom[6872] = 8'hea ;
            rom[6873] = 8'hf5 ;
            rom[6874] = 8'he0 ;
            rom[6875] = 8'h14 ;
            rom[6876] = 8'h04 ;
            rom[6877] = 8'h18 ;
            rom[6878] = 8'h1c ;
            rom[6879] = 8'h1b ;
            rom[6880] = 8'h02 ;
            rom[6881] = 8'hf6 ;
            rom[6882] = 8'h0d ;
            rom[6883] = 8'h00 ;
            rom[6884] = 8'h03 ;
            rom[6885] = 8'h20 ;
            rom[6886] = 8'he4 ;
            rom[6887] = 8'he3 ;
            rom[6888] = 8'he6 ;
            rom[6889] = 8'hf7 ;
            rom[6890] = 8'h0d ;
            rom[6891] = 8'hed ;
            rom[6892] = 8'h2a ;
            rom[6893] = 8'h19 ;
            rom[6894] = 8'hd4 ;
            rom[6895] = 8'h29 ;
            rom[6896] = 8'hfe ;
            rom[6897] = 8'h0a ;
            rom[6898] = 8'hf4 ;
            rom[6899] = 8'hff ;
            rom[6900] = 8'h12 ;
            rom[6901] = 8'h00 ;
            rom[6902] = 8'h13 ;
            rom[6903] = 8'hff ;
            rom[6904] = 8'hff ;
            rom[6905] = 8'h09 ;
            rom[6906] = 8'h0e ;
            rom[6907] = 8'hfc ;
            rom[6908] = 8'h0d ;
            rom[6909] = 8'h29 ;
            rom[6910] = 8'hf8 ;
            rom[6911] = 8'h07 ;
            rom[6912] = 8'hf5 ;
            rom[6913] = 8'hf5 ;
            rom[6914] = 8'hf9 ;
            rom[6915] = 8'hf2 ;
            rom[6916] = 8'h2d ;
            rom[6917] = 8'h17 ;
            rom[6918] = 8'hd2 ;
            rom[6919] = 8'hf9 ;
            rom[6920] = 8'hc2 ;
            rom[6921] = 8'h1a ;
            rom[6922] = 8'hfa ;
            rom[6923] = 8'hfd ;
            rom[6924] = 8'h0c ;
            rom[6925] = 8'hf3 ;
            rom[6926] = 8'h00 ;
            rom[6927] = 8'hf6 ;
            rom[6928] = 8'hf9 ;
            rom[6929] = 8'hf8 ;
            rom[6930] = 8'hde ;
            rom[6931] = 8'h04 ;
            rom[6932] = 8'h05 ;
            rom[6933] = 8'h16 ;
            rom[6934] = 8'h0a ;
            rom[6935] = 8'hf8 ;
            rom[6936] = 8'hf3 ;
            rom[6937] = 8'he8 ;
            rom[6938] = 8'hf2 ;
            rom[6939] = 8'hff ;
            rom[6940] = 8'hc9 ;
            rom[6941] = 8'he7 ;
            rom[6942] = 8'h03 ;
            rom[6943] = 8'h11 ;
            rom[6944] = 8'he8 ;
            rom[6945] = 8'he1 ;
            rom[6946] = 8'hfd ;
            rom[6947] = 8'h06 ;
            rom[6948] = 8'h05 ;
            rom[6949] = 8'h18 ;
            rom[6950] = 8'he0 ;
            rom[6951] = 8'h1c ;
            rom[6952] = 8'h11 ;
            rom[6953] = 8'hfb ;
            rom[6954] = 8'hf4 ;
            rom[6955] = 8'h0a ;
            rom[6956] = 8'hfe ;
            rom[6957] = 8'h23 ;
            rom[6958] = 8'he9 ;
            rom[6959] = 8'h18 ;
            rom[6960] = 8'hff ;
            rom[6961] = 8'hf6 ;
            rom[6962] = 8'hfe ;
            rom[6963] = 8'hed ;
            rom[6964] = 8'h07 ;
            rom[6965] = 8'hdf ;
            rom[6966] = 8'h1e ;
            rom[6967] = 8'h06 ;
            rom[6968] = 8'h01 ;
            rom[6969] = 8'he6 ;
            rom[6970] = 8'he5 ;
            rom[6971] = 8'h09 ;
            rom[6972] = 8'hc1 ;
            rom[6973] = 8'hf5 ;
            rom[6974] = 8'h17 ;
            rom[6975] = 8'h22 ;
            rom[6976] = 8'h09 ;
            rom[6977] = 8'h17 ;
            rom[6978] = 8'h15 ;
            rom[6979] = 8'hfb ;
            rom[6980] = 8'he3 ;
            rom[6981] = 8'h08 ;
            rom[6982] = 8'hf3 ;
            rom[6983] = 8'he2 ;
            rom[6984] = 8'he7 ;
            rom[6985] = 8'he8 ;
            rom[6986] = 8'h14 ;
            rom[6987] = 8'hff ;
            rom[6988] = 8'hd6 ;
            rom[6989] = 8'hfa ;
            rom[6990] = 8'h09 ;
            rom[6991] = 8'h11 ;
            rom[6992] = 8'hfb ;
            rom[6993] = 8'he7 ;
            rom[6994] = 8'h03 ;
            rom[6995] = 8'hc4 ;
            rom[6996] = 8'hda ;
            rom[6997] = 8'h02 ;
            rom[6998] = 8'h0f ;
            rom[6999] = 8'h05 ;
            rom[7000] = 8'hee ;
            rom[7001] = 8'h01 ;
            rom[7002] = 8'hee ;
            rom[7003] = 8'hf6 ;
            rom[7004] = 8'hef ;
            rom[7005] = 8'h16 ;
            rom[7006] = 8'h0f ;
            rom[7007] = 8'h02 ;
            rom[7008] = 8'h03 ;
            rom[7009] = 8'hfb ;
            rom[7010] = 8'h0b ;
            rom[7011] = 8'h1e ;
            rom[7012] = 8'he2 ;
            rom[7013] = 8'h01 ;
            rom[7014] = 8'h05 ;
            rom[7015] = 8'h15 ;
            rom[7016] = 8'hf3 ;
            rom[7017] = 8'hff ;
            rom[7018] = 8'hfd ;
            rom[7019] = 8'hf3 ;
            rom[7020] = 8'hde ;
            rom[7021] = 8'h1b ;
            rom[7022] = 8'h05 ;
            rom[7023] = 8'hd1 ;
            rom[7024] = 8'h09 ;
            rom[7025] = 8'h10 ;
            rom[7026] = 8'h0a ;
            rom[7027] = 8'hed ;
            rom[7028] = 8'he4 ;
            rom[7029] = 8'he7 ;
            rom[7030] = 8'hfc ;
            rom[7031] = 8'h21 ;
            rom[7032] = 8'h0f ;
            rom[7033] = 8'hfd ;
            rom[7034] = 8'hf7 ;
            rom[7035] = 8'hf8 ;
            rom[7036] = 8'hfe ;
            rom[7037] = 8'h0c ;
            rom[7038] = 8'hf5 ;
            rom[7039] = 8'h01 ;
            rom[7040] = 8'h31 ;
            rom[7041] = 8'h23 ;
            rom[7042] = 8'he7 ;
            rom[7043] = 8'h03 ;
            rom[7044] = 8'hef ;
            rom[7045] = 8'h2a ;
            rom[7046] = 8'hfa ;
            rom[7047] = 8'hed ;
            rom[7048] = 8'he8 ;
            rom[7049] = 8'hef ;
            rom[7050] = 8'h01 ;
            rom[7051] = 8'h07 ;
            rom[7052] = 8'hfd ;
            rom[7053] = 8'hf8 ;
            rom[7054] = 8'h1d ;
            rom[7055] = 8'he7 ;
            rom[7056] = 8'hf4 ;
            rom[7057] = 8'hed ;
            rom[7058] = 8'h03 ;
            rom[7059] = 8'hd6 ;
            rom[7060] = 8'hfa ;
            rom[7061] = 8'h1c ;
            rom[7062] = 8'hf7 ;
            rom[7063] = 8'ha9 ;
            rom[7064] = 8'hd7 ;
            rom[7065] = 8'h0e ;
            rom[7066] = 8'hf8 ;
            rom[7067] = 8'hf3 ;
            rom[7068] = 8'he2 ;
            rom[7069] = 8'h08 ;
            rom[7070] = 8'hf4 ;
            rom[7071] = 8'h00 ;
            rom[7072] = 8'h0c ;
            rom[7073] = 8'h08 ;
            rom[7074] = 8'h12 ;
            rom[7075] = 8'h3b ;
            rom[7076] = 8'h11 ;
            rom[7077] = 8'h1b ;
            rom[7078] = 8'hde ;
            rom[7079] = 8'h0d ;
            rom[7080] = 8'h0f ;
            rom[7081] = 8'hfe ;
            rom[7082] = 8'hf3 ;
            rom[7083] = 8'h1c ;
            rom[7084] = 8'hee ;
            rom[7085] = 8'h1b ;
            rom[7086] = 8'h1e ;
            rom[7087] = 8'hcf ;
            rom[7088] = 8'h24 ;
            rom[7089] = 8'h11 ;
            rom[7090] = 8'hf7 ;
            rom[7091] = 8'h10 ;
            rom[7092] = 8'h03 ;
            rom[7093] = 8'hdc ;
            rom[7094] = 8'hfb ;
            rom[7095] = 8'hf7 ;
            rom[7096] = 8'h00 ;
            rom[7097] = 8'h08 ;
            rom[7098] = 8'h15 ;
            rom[7099] = 8'h0b ;
            rom[7100] = 8'h13 ;
            rom[7101] = 8'hde ;
            rom[7102] = 8'h0d ;
            rom[7103] = 8'hec ;
            rom[7104] = 8'hff ;
            rom[7105] = 8'h00 ;
            rom[7106] = 8'hf6 ;
            rom[7107] = 8'h08 ;
            rom[7108] = 8'h21 ;
            rom[7109] = 8'h0e ;
            rom[7110] = 8'hf1 ;
            rom[7111] = 8'hfd ;
            rom[7112] = 8'hde ;
            rom[7113] = 8'h1a ;
            rom[7114] = 8'hf8 ;
            rom[7115] = 8'h10 ;
            rom[7116] = 8'h12 ;
            rom[7117] = 8'h13 ;
            rom[7118] = 8'h0b ;
            rom[7119] = 8'hf0 ;
            rom[7120] = 8'h03 ;
            rom[7121] = 8'hc5 ;
            rom[7122] = 8'he6 ;
            rom[7123] = 8'hd8 ;
            rom[7124] = 8'hf9 ;
            rom[7125] = 8'hff ;
            rom[7126] = 8'h1c ;
            rom[7127] = 8'hec ;
            rom[7128] = 8'hdb ;
            rom[7129] = 8'h11 ;
            rom[7130] = 8'he1 ;
            rom[7131] = 8'h0f ;
            rom[7132] = 8'hfe ;
            rom[7133] = 8'hf9 ;
            rom[7134] = 8'h0e ;
            rom[7135] = 8'h01 ;
            rom[7136] = 8'hf0 ;
            rom[7137] = 8'h06 ;
            rom[7138] = 8'h03 ;
            rom[7139] = 8'hff ;
            rom[7140] = 8'hd8 ;
            rom[7141] = 8'h08 ;
            rom[7142] = 8'he0 ;
            rom[7143] = 8'he3 ;
            rom[7144] = 8'hfc ;
            rom[7145] = 8'h01 ;
            rom[7146] = 8'h00 ;
            rom[7147] = 8'h06 ;
            rom[7148] = 8'hf0 ;
            rom[7149] = 8'h32 ;
            rom[7150] = 8'h04 ;
            rom[7151] = 8'h15 ;
            rom[7152] = 8'hed ;
            rom[7153] = 8'h02 ;
            rom[7154] = 8'hf3 ;
            rom[7155] = 8'h0a ;
            rom[7156] = 8'hf1 ;
            rom[7157] = 8'hf2 ;
            rom[7158] = 8'h0a ;
            rom[7159] = 8'h01 ;
            rom[7160] = 8'hef ;
            rom[7161] = 8'hf6 ;
            rom[7162] = 8'hfa ;
            rom[7163] = 8'h04 ;
            rom[7164] = 8'he0 ;
            rom[7165] = 8'h1f ;
            rom[7166] = 8'h06 ;
            rom[7167] = 8'h09 ;
            rom[7168] = 8'hfb ;
            rom[7169] = 8'h0d ;
            rom[7170] = 8'hd6 ;
            rom[7171] = 8'h1b ;
            rom[7172] = 8'h29 ;
            rom[7173] = 8'hf0 ;
            rom[7174] = 8'hfb ;
            rom[7175] = 8'h11 ;
            rom[7176] = 8'hf5 ;
            rom[7177] = 8'h02 ;
            rom[7178] = 8'hef ;
            rom[7179] = 8'h00 ;
            rom[7180] = 8'hf9 ;
            rom[7181] = 8'h19 ;
            rom[7182] = 8'he6 ;
            rom[7183] = 8'h03 ;
            rom[7184] = 8'hf6 ;
            rom[7185] = 8'h08 ;
            rom[7186] = 8'h25 ;
            rom[7187] = 8'hfd ;
            rom[7188] = 8'h0d ;
            rom[7189] = 8'hfd ;
            rom[7190] = 8'he4 ;
            rom[7191] = 8'hf9 ;
            rom[7192] = 8'h06 ;
            rom[7193] = 8'hf7 ;
            rom[7194] = 8'hff ;
            rom[7195] = 8'hff ;
            rom[7196] = 8'hf7 ;
            rom[7197] = 8'hed ;
            rom[7198] = 8'h02 ;
            rom[7199] = 8'h17 ;
            rom[7200] = 8'he5 ;
            rom[7201] = 8'h0d ;
            rom[7202] = 8'h06 ;
            rom[7203] = 8'hfd ;
            rom[7204] = 8'hf3 ;
            rom[7205] = 8'h0a ;
            rom[7206] = 8'h05 ;
            rom[7207] = 8'hfc ;
            rom[7208] = 8'hf2 ;
            rom[7209] = 8'h08 ;
            rom[7210] = 8'hfe ;
            rom[7211] = 8'hf0 ;
            rom[7212] = 8'heb ;
            rom[7213] = 8'h08 ;
            rom[7214] = 8'hea ;
            rom[7215] = 8'h12 ;
            rom[7216] = 8'h17 ;
            rom[7217] = 8'h08 ;
            rom[7218] = 8'hdc ;
            rom[7219] = 8'h09 ;
            rom[7220] = 8'h0d ;
            rom[7221] = 8'ha1 ;
            rom[7222] = 8'hfe ;
            rom[7223] = 8'hf9 ;
            rom[7224] = 8'hd5 ;
            rom[7225] = 8'he9 ;
            rom[7226] = 8'hf0 ;
            rom[7227] = 8'h33 ;
            rom[7228] = 8'hc9 ;
            rom[7229] = 8'he2 ;
            rom[7230] = 8'h15 ;
            rom[7231] = 8'h18 ;
            rom[7232] = 8'h0d ;
            rom[7233] = 8'hfa ;
            rom[7234] = 8'h1c ;
            rom[7235] = 8'h01 ;
            rom[7236] = 8'h0b ;
            rom[7237] = 8'h03 ;
            rom[7238] = 8'h1f ;
            rom[7239] = 8'h14 ;
            rom[7240] = 8'hf2 ;
            rom[7241] = 8'hf9 ;
            rom[7242] = 8'h02 ;
            rom[7243] = 8'hd6 ;
            rom[7244] = 8'h00 ;
            rom[7245] = 8'hf6 ;
            rom[7246] = 8'hf4 ;
            rom[7247] = 8'h08 ;
            rom[7248] = 8'hf2 ;
            rom[7249] = 8'h0f ;
            rom[7250] = 8'hf8 ;
            rom[7251] = 8'h24 ;
            rom[7252] = 8'h02 ;
            rom[7253] = 8'h18 ;
            rom[7254] = 8'h05 ;
            rom[7255] = 8'h12 ;
            rom[7256] = 8'h0a ;
            rom[7257] = 8'h08 ;
            rom[7258] = 8'hf0 ;
            rom[7259] = 8'h00 ;
            rom[7260] = 8'hef ;
            rom[7261] = 8'h2d ;
            rom[7262] = 8'h12 ;
            rom[7263] = 8'h0c ;
            rom[7264] = 8'hed ;
            rom[7265] = 8'hf8 ;
            rom[7266] = 8'hde ;
            rom[7267] = 8'h04 ;
            rom[7268] = 8'h23 ;
            rom[7269] = 8'h2c ;
            rom[7270] = 8'h2b ;
            rom[7271] = 8'he5 ;
            rom[7272] = 8'h0f ;
            rom[7273] = 8'hec ;
            rom[7274] = 8'hfb ;
            rom[7275] = 8'h05 ;
            rom[7276] = 8'h0e ;
            rom[7277] = 8'h0e ;
            rom[7278] = 8'h02 ;
            rom[7279] = 8'h02 ;
            rom[7280] = 8'h2d ;
            rom[7281] = 8'h07 ;
            rom[7282] = 8'h20 ;
            rom[7283] = 8'hee ;
            rom[7284] = 8'h2b ;
            rom[7285] = 8'h00 ;
            rom[7286] = 8'hff ;
            rom[7287] = 8'h12 ;
            rom[7288] = 8'h0a ;
            rom[7289] = 8'hf4 ;
            rom[7290] = 8'hef ;
            rom[7291] = 8'h13 ;
            rom[7292] = 8'hee ;
            rom[7293] = 8'hf6 ;
            rom[7294] = 8'h05 ;
            rom[7295] = 8'hf4 ;
            rom[7296] = 8'h07 ;
            rom[7297] = 8'hf6 ;
            rom[7298] = 8'hee ;
            rom[7299] = 8'hee ;
            rom[7300] = 8'h0c ;
            rom[7301] = 8'h26 ;
            rom[7302] = 8'h13 ;
            rom[7303] = 8'h09 ;
            rom[7304] = 8'hca ;
            rom[7305] = 8'h0c ;
            rom[7306] = 8'h08 ;
            rom[7307] = 8'h13 ;
            rom[7308] = 8'hfa ;
            rom[7309] = 8'hcd ;
            rom[7310] = 8'h27 ;
            rom[7311] = 8'hf5 ;
            rom[7312] = 8'hf8 ;
            rom[7313] = 8'hf5 ;
            rom[7314] = 8'hf5 ;
            rom[7315] = 8'h1c ;
            rom[7316] = 8'hff ;
            rom[7317] = 8'h10 ;
            rom[7318] = 8'hfb ;
            rom[7319] = 8'hf6 ;
            rom[7320] = 8'hf1 ;
            rom[7321] = 8'h01 ;
            rom[7322] = 8'h0f ;
            rom[7323] = 8'h1c ;
            rom[7324] = 8'hde ;
            rom[7325] = 8'h06 ;
            rom[7326] = 8'hf6 ;
            rom[7327] = 8'hfc ;
            rom[7328] = 8'he6 ;
            rom[7329] = 8'hff ;
            rom[7330] = 8'hf2 ;
            rom[7331] = 8'h13 ;
            rom[7332] = 8'h16 ;
            rom[7333] = 8'h17 ;
            rom[7334] = 8'h12 ;
            rom[7335] = 8'h1c ;
            rom[7336] = 8'h0f ;
            rom[7337] = 8'hf9 ;
            rom[7338] = 8'h05 ;
            rom[7339] = 8'h11 ;
            rom[7340] = 8'he7 ;
            rom[7341] = 8'hff ;
            rom[7342] = 8'h00 ;
            rom[7343] = 8'hdf ;
            rom[7344] = 8'hf4 ;
            rom[7345] = 8'h18 ;
            rom[7346] = 8'h02 ;
            rom[7347] = 8'h0c ;
            rom[7348] = 8'h04 ;
            rom[7349] = 8'hdb ;
            rom[7350] = 8'h18 ;
            rom[7351] = 8'h10 ;
            rom[7352] = 8'hf2 ;
            rom[7353] = 8'he9 ;
            rom[7354] = 8'h16 ;
            rom[7355] = 8'h12 ;
            rom[7356] = 8'hd6 ;
            rom[7357] = 8'hf3 ;
            rom[7358] = 8'hef ;
            rom[7359] = 8'hf3 ;
            rom[7360] = 8'he9 ;
            rom[7361] = 8'h19 ;
            rom[7362] = 8'hef ;
            rom[7363] = 8'hfc ;
            rom[7364] = 8'hf9 ;
            rom[7365] = 8'hea ;
            rom[7366] = 8'h0b ;
            rom[7367] = 8'hf6 ;
            rom[7368] = 8'hf7 ;
            rom[7369] = 8'hdf ;
            rom[7370] = 8'hbc ;
            rom[7371] = 8'hf3 ;
            rom[7372] = 8'he6 ;
            rom[7373] = 8'hff ;
            rom[7374] = 8'hf7 ;
            rom[7375] = 8'hfd ;
            rom[7376] = 8'h15 ;
            rom[7377] = 8'hf6 ;
            rom[7378] = 8'he7 ;
            rom[7379] = 8'h00 ;
            rom[7380] = 8'hde ;
            rom[7381] = 8'h0a ;
            rom[7382] = 8'hff ;
            rom[7383] = 8'hf4 ;
            rom[7384] = 8'hf8 ;
            rom[7385] = 8'hf9 ;
            rom[7386] = 8'hf0 ;
            rom[7387] = 8'h02 ;
            rom[7388] = 8'he1 ;
            rom[7389] = 8'hf9 ;
            rom[7390] = 8'h20 ;
            rom[7391] = 8'h1a ;
            rom[7392] = 8'h00 ;
            rom[7393] = 8'hfe ;
            rom[7394] = 8'hfa ;
            rom[7395] = 8'h00 ;
            rom[7396] = 8'hf6 ;
            rom[7397] = 8'h12 ;
            rom[7398] = 8'hf2 ;
            rom[7399] = 8'h09 ;
            rom[7400] = 8'hfe ;
            rom[7401] = 8'h02 ;
            rom[7402] = 8'he3 ;
            rom[7403] = 8'hf0 ;
            rom[7404] = 8'hdf ;
            rom[7405] = 8'h03 ;
            rom[7406] = 8'hbd ;
            rom[7407] = 8'h0c ;
            rom[7408] = 8'h1f ;
            rom[7409] = 8'hed ;
            rom[7410] = 8'h03 ;
            rom[7411] = 8'hfb ;
            rom[7412] = 8'h03 ;
            rom[7413] = 8'hf8 ;
            rom[7414] = 8'hce ;
            rom[7415] = 8'h10 ;
            rom[7416] = 8'hf8 ;
            rom[7417] = 8'h08 ;
            rom[7418] = 8'hef ;
            rom[7419] = 8'hfa ;
            rom[7420] = 8'h15 ;
            rom[7421] = 8'h12 ;
            rom[7422] = 8'hfb ;
            rom[7423] = 8'h01 ;
            rom[7424] = 8'h31 ;
            rom[7425] = 8'h0d ;
            rom[7426] = 8'h04 ;
            rom[7427] = 8'he4 ;
            rom[7428] = 8'h1a ;
            rom[7429] = 8'h05 ;
            rom[7430] = 8'hfa ;
            rom[7431] = 8'heb ;
            rom[7432] = 8'he7 ;
            rom[7433] = 8'hfb ;
            rom[7434] = 8'hfa ;
            rom[7435] = 8'he4 ;
            rom[7436] = 8'h02 ;
            rom[7437] = 8'hf1 ;
            rom[7438] = 8'hd6 ;
            rom[7439] = 8'h06 ;
            rom[7440] = 8'h09 ;
            rom[7441] = 8'hfb ;
            rom[7442] = 8'h2c ;
            rom[7443] = 8'h1a ;
            rom[7444] = 8'he9 ;
            rom[7445] = 8'hfa ;
            rom[7446] = 8'hf1 ;
            rom[7447] = 8'hf9 ;
            rom[7448] = 8'hfa ;
            rom[7449] = 8'hd3 ;
            rom[7450] = 8'hf1 ;
            rom[7451] = 8'hf6 ;
            rom[7452] = 8'h06 ;
            rom[7453] = 8'hfd ;
            rom[7454] = 8'hd6 ;
            rom[7455] = 8'h02 ;
            rom[7456] = 8'hfc ;
            rom[7457] = 8'h1b ;
            rom[7458] = 8'h18 ;
            rom[7459] = 8'hf4 ;
            rom[7460] = 8'h23 ;
            rom[7461] = 8'h12 ;
            rom[7462] = 8'h09 ;
            rom[7463] = 8'h02 ;
            rom[7464] = 8'h12 ;
            rom[7465] = 8'hf0 ;
            rom[7466] = 8'hfe ;
            rom[7467] = 8'hef ;
            rom[7468] = 8'hea ;
            rom[7469] = 8'h05 ;
            rom[7470] = 8'h02 ;
            rom[7471] = 8'hf6 ;
            rom[7472] = 8'h0c ;
            rom[7473] = 8'h09 ;
            rom[7474] = 8'h1a ;
            rom[7475] = 8'hff ;
            rom[7476] = 8'h07 ;
            rom[7477] = 8'hda ;
            rom[7478] = 8'h09 ;
            rom[7479] = 8'h0d ;
            rom[7480] = 8'hf5 ;
            rom[7481] = 8'hb9 ;
            rom[7482] = 8'he1 ;
            rom[7483] = 8'h19 ;
            rom[7484] = 8'h0c ;
            rom[7485] = 8'hdf ;
            rom[7486] = 8'hfd ;
            rom[7487] = 8'hf0 ;
            rom[7488] = 8'h13 ;
            rom[7489] = 8'hfc ;
            rom[7490] = 8'he4 ;
            rom[7491] = 8'h16 ;
            rom[7492] = 8'h28 ;
            rom[7493] = 8'hcd ;
            rom[7494] = 8'h18 ;
            rom[7495] = 8'h03 ;
            rom[7496] = 8'h13 ;
            rom[7497] = 8'hda ;
            rom[7498] = 8'hf1 ;
            rom[7499] = 8'h05 ;
            rom[7500] = 8'h0a ;
            rom[7501] = 8'h01 ;
            rom[7502] = 8'h00 ;
            rom[7503] = 8'he7 ;
            rom[7504] = 8'h23 ;
            rom[7505] = 8'h0d ;
            rom[7506] = 8'h07 ;
            rom[7507] = 8'h01 ;
            rom[7508] = 8'h1c ;
            rom[7509] = 8'hfb ;
            rom[7510] = 8'hf8 ;
            rom[7511] = 8'h07 ;
            rom[7512] = 8'hfd ;
            rom[7513] = 8'he8 ;
            rom[7514] = 8'h0d ;
            rom[7515] = 8'h06 ;
            rom[7516] = 8'he8 ;
            rom[7517] = 8'hfa ;
            rom[7518] = 8'h1e ;
            rom[7519] = 8'h19 ;
            rom[7520] = 8'he3 ;
            rom[7521] = 8'hee ;
            rom[7522] = 8'hd4 ;
            rom[7523] = 8'hf9 ;
            rom[7524] = 8'hdb ;
            rom[7525] = 8'hfe ;
            rom[7526] = 8'hc0 ;
            rom[7527] = 8'hfe ;
            rom[7528] = 8'hf5 ;
            rom[7529] = 8'hef ;
            rom[7530] = 8'h1d ;
            rom[7531] = 8'h01 ;
            rom[7532] = 8'hfb ;
            rom[7533] = 8'h06 ;
            rom[7534] = 8'he8 ;
            rom[7535] = 8'h1f ;
            rom[7536] = 8'h0d ;
            rom[7537] = 8'h1b ;
            rom[7538] = 8'he4 ;
            rom[7539] = 8'hf9 ;
            rom[7540] = 8'hdf ;
            rom[7541] = 8'hf2 ;
            rom[7542] = 8'h07 ;
            rom[7543] = 8'h0a ;
            rom[7544] = 8'hd2 ;
            rom[7545] = 8'he5 ;
            rom[7546] = 8'h08 ;
            rom[7547] = 8'h2d ;
            rom[7548] = 8'h08 ;
            rom[7549] = 8'hff ;
            rom[7550] = 8'h18 ;
            rom[7551] = 8'hfe ;
            rom[7552] = 8'h08 ;
            rom[7553] = 8'hfd ;
            rom[7554] = 8'hfe ;
            rom[7555] = 8'h0d ;
            rom[7556] = 8'h19 ;
            rom[7557] = 8'h1b ;
            rom[7558] = 8'hfb ;
            rom[7559] = 8'he4 ;
            rom[7560] = 8'h0c ;
            rom[7561] = 8'he8 ;
            rom[7562] = 8'h18 ;
            rom[7563] = 8'hf3 ;
            rom[7564] = 8'h21 ;
            rom[7565] = 8'hfb ;
            rom[7566] = 8'he8 ;
            rom[7567] = 8'hf6 ;
            rom[7568] = 8'hf9 ;
            rom[7569] = 8'h14 ;
            rom[7570] = 8'hec ;
            rom[7571] = 8'hec ;
            rom[7572] = 8'h0a ;
            rom[7573] = 8'hf1 ;
            rom[7574] = 8'hf5 ;
            rom[7575] = 8'h18 ;
            rom[7576] = 8'h09 ;
            rom[7577] = 8'hcd ;
            rom[7578] = 8'hd9 ;
            rom[7579] = 8'h15 ;
            rom[7580] = 8'h05 ;
            rom[7581] = 8'h11 ;
            rom[7582] = 8'hfd ;
            rom[7583] = 8'h17 ;
            rom[7584] = 8'hf3 ;
            rom[7585] = 8'hfe ;
            rom[7586] = 8'hcc ;
            rom[7587] = 8'h09 ;
            rom[7588] = 8'h16 ;
            rom[7589] = 8'he5 ;
            rom[7590] = 8'hfa ;
            rom[7591] = 8'h26 ;
            rom[7592] = 8'hfc ;
            rom[7593] = 8'hf4 ;
            rom[7594] = 8'h04 ;
            rom[7595] = 8'hfe ;
            rom[7596] = 8'hf3 ;
            rom[7597] = 8'h01 ;
            rom[7598] = 8'h0e ;
            rom[7599] = 8'hea ;
            rom[7600] = 8'hf5 ;
            rom[7601] = 8'hf4 ;
            rom[7602] = 8'hea ;
            rom[7603] = 8'hff ;
            rom[7604] = 8'hcb ;
            rom[7605] = 8'h02 ;
            rom[7606] = 8'h1f ;
            rom[7607] = 8'h1b ;
            rom[7608] = 8'h0e ;
            rom[7609] = 8'h0b ;
            rom[7610] = 8'hfc ;
            rom[7611] = 8'h02 ;
            rom[7612] = 8'h09 ;
            rom[7613] = 8'hdb ;
            rom[7614] = 8'h15 ;
            rom[7615] = 8'hf8 ;
            rom[7616] = 8'hf3 ;
            rom[7617] = 8'h1d ;
            rom[7618] = 8'he6 ;
            rom[7619] = 8'h07 ;
            rom[7620] = 8'h10 ;
            rom[7621] = 8'hfa ;
            rom[7622] = 8'h0c ;
            rom[7623] = 8'h0b ;
            rom[7624] = 8'h0c ;
            rom[7625] = 8'hf4 ;
            rom[7626] = 8'hd0 ;
            rom[7627] = 8'h11 ;
            rom[7628] = 8'hed ;
            rom[7629] = 8'hf2 ;
            rom[7630] = 8'h14 ;
            rom[7631] = 8'hf0 ;
            rom[7632] = 8'h19 ;
            rom[7633] = 8'h13 ;
            rom[7634] = 8'h15 ;
            rom[7635] = 8'h0c ;
            rom[7636] = 8'h05 ;
            rom[7637] = 8'h03 ;
            rom[7638] = 8'hfd ;
            rom[7639] = 8'h25 ;
            rom[7640] = 8'he7 ;
            rom[7641] = 8'h00 ;
            rom[7642] = 8'hf4 ;
            rom[7643] = 8'hf8 ;
            rom[7644] = 8'hdb ;
            rom[7645] = 8'h09 ;
            rom[7646] = 8'h08 ;
            rom[7647] = 8'h0d ;
            rom[7648] = 8'he2 ;
            rom[7649] = 8'he4 ;
            rom[7650] = 8'heb ;
            rom[7651] = 8'h01 ;
            rom[7652] = 8'h04 ;
            rom[7653] = 8'hec ;
            rom[7654] = 8'hd5 ;
            rom[7655] = 8'hed ;
            rom[7656] = 8'h02 ;
            rom[7657] = 8'hf5 ;
            rom[7658] = 8'hfe ;
            rom[7659] = 8'h0c ;
            rom[7660] = 8'hef ;
            rom[7661] = 8'hea ;
            rom[7662] = 8'hf3 ;
            rom[7663] = 8'h16 ;
            rom[7664] = 8'hfa ;
            rom[7665] = 8'h1f ;
            rom[7666] = 8'h0f ;
            rom[7667] = 8'h02 ;
            rom[7668] = 8'he2 ;
            rom[7669] = 8'h06 ;
            rom[7670] = 8'h06 ;
            rom[7671] = 8'h02 ;
            rom[7672] = 8'hb3 ;
            rom[7673] = 8'hfd ;
            rom[7674] = 8'h21 ;
            rom[7675] = 8'h41 ;
            rom[7676] = 8'he2 ;
            rom[7677] = 8'hf9 ;
            rom[7678] = 8'hf6 ;
            rom[7679] = 8'h23 ;
            rom[7680] = 8'hf7 ;
            rom[7681] = 8'hd6 ;
            rom[7682] = 8'h13 ;
            rom[7683] = 8'hf0 ;
            rom[7684] = 8'h0c ;
            rom[7685] = 8'h1a ;
            rom[7686] = 8'hdd ;
            rom[7687] = 8'hf0 ;
            rom[7688] = 8'hd2 ;
            rom[7689] = 8'hf1 ;
            rom[7690] = 8'h04 ;
            rom[7691] = 8'heb ;
            rom[7692] = 8'h16 ;
            rom[7693] = 8'he0 ;
            rom[7694] = 8'hf5 ;
            rom[7695] = 8'hd7 ;
            rom[7696] = 8'h02 ;
            rom[7697] = 8'h02 ;
            rom[7698] = 8'hd8 ;
            rom[7699] = 8'h04 ;
            rom[7700] = 8'hed ;
            rom[7701] = 8'h11 ;
            rom[7702] = 8'hfc ;
            rom[7703] = 8'hf7 ;
            rom[7704] = 8'h17 ;
            rom[7705] = 8'hf6 ;
            rom[7706] = 8'he7 ;
            rom[7707] = 8'hea ;
            rom[7708] = 8'h13 ;
            rom[7709] = 8'h14 ;
            rom[7710] = 8'h02 ;
            rom[7711] = 8'hdc ;
            rom[7712] = 8'h05 ;
            rom[7713] = 8'hf2 ;
            rom[7714] = 8'hca ;
            rom[7715] = 8'h22 ;
            rom[7716] = 8'hed ;
            rom[7717] = 8'h0b ;
            rom[7718] = 8'h18 ;
            rom[7719] = 8'h1d ;
            rom[7720] = 8'h1f ;
            rom[7721] = 8'hc4 ;
            rom[7722] = 8'h06 ;
            rom[7723] = 8'h0e ;
            rom[7724] = 8'hff ;
            rom[7725] = 8'h13 ;
            rom[7726] = 8'h0e ;
            rom[7727] = 8'h12 ;
            rom[7728] = 8'h03 ;
            rom[7729] = 8'h01 ;
            rom[7730] = 8'h28 ;
            rom[7731] = 8'hf3 ;
            rom[7732] = 8'he9 ;
            rom[7733] = 8'hed ;
            rom[7734] = 8'hf7 ;
            rom[7735] = 8'h13 ;
            rom[7736] = 8'h05 ;
            rom[7737] = 8'hcc ;
            rom[7738] = 8'hf7 ;
            rom[7739] = 8'h17 ;
            rom[7740] = 8'hf9 ;
            rom[7741] = 8'hd1 ;
            rom[7742] = 8'h1b ;
            rom[7743] = 8'hf0 ;
            rom[7744] = 8'hee ;
            rom[7745] = 8'h0f ;
            rom[7746] = 8'hf6 ;
            rom[7747] = 8'h1c ;
            rom[7748] = 8'h08 ;
            rom[7749] = 8'heb ;
            rom[7750] = 8'h0f ;
            rom[7751] = 8'h0d ;
            rom[7752] = 8'he6 ;
            rom[7753] = 8'hbf ;
            rom[7754] = 8'hbd ;
            rom[7755] = 8'hf9 ;
            rom[7756] = 8'he8 ;
            rom[7757] = 8'he7 ;
            rom[7758] = 8'h03 ;
            rom[7759] = 8'hfb ;
            rom[7760] = 8'hf1 ;
            rom[7761] = 8'h0a ;
            rom[7762] = 8'hff ;
            rom[7763] = 8'hf4 ;
            rom[7764] = 8'hed ;
            rom[7765] = 8'h18 ;
            rom[7766] = 8'he8 ;
            rom[7767] = 8'hff ;
            rom[7768] = 8'h19 ;
            rom[7769] = 8'hd6 ;
            rom[7770] = 8'h0e ;
            rom[7771] = 8'hfd ;
            rom[7772] = 8'he4 ;
            rom[7773] = 8'h1e ;
            rom[7774] = 8'hf9 ;
            rom[7775] = 8'hde ;
            rom[7776] = 8'h12 ;
            rom[7777] = 8'he7 ;
            rom[7778] = 8'hf1 ;
            rom[7779] = 8'hed ;
            rom[7780] = 8'hea ;
            rom[7781] = 8'h10 ;
            rom[7782] = 8'hf4 ;
            rom[7783] = 8'h00 ;
            rom[7784] = 8'h15 ;
            rom[7785] = 8'hb3 ;
            rom[7786] = 8'hc9 ;
            rom[7787] = 8'h01 ;
            rom[7788] = 8'hf5 ;
            rom[7789] = 8'h01 ;
            rom[7790] = 8'hdb ;
            rom[7791] = 8'hff ;
            rom[7792] = 8'h05 ;
            rom[7793] = 8'he2 ;
            rom[7794] = 8'h0b ;
            rom[7795] = 8'hf9 ;
            rom[7796] = 8'hd8 ;
            rom[7797] = 8'h11 ;
            rom[7798] = 8'hce ;
            rom[7799] = 8'h08 ;
            rom[7800] = 8'hf7 ;
            rom[7801] = 8'h03 ;
            rom[7802] = 8'h0c ;
            rom[7803] = 8'h0c ;
            rom[7804] = 8'h0a ;
            rom[7805] = 8'h0b ;
            rom[7806] = 8'h12 ;
            rom[7807] = 8'hf8 ;
            rom[7808] = 8'hea ;
            rom[7809] = 8'h0b ;
            rom[7810] = 8'heb ;
            rom[7811] = 8'h12 ;
            rom[7812] = 8'h1c ;
            rom[7813] = 8'heb ;
            rom[7814] = 8'h0e ;
            rom[7815] = 8'hfe ;
            rom[7816] = 8'hfa ;
            rom[7817] = 8'ha2 ;
            rom[7818] = 8'hd6 ;
            rom[7819] = 8'hed ;
            rom[7820] = 8'h0e ;
            rom[7821] = 8'hf0 ;
            rom[7822] = 8'h13 ;
            rom[7823] = 8'hf6 ;
            rom[7824] = 8'hf0 ;
            rom[7825] = 8'h12 ;
            rom[7826] = 8'h07 ;
            rom[7827] = 8'hd6 ;
            rom[7828] = 8'hfe ;
            rom[7829] = 8'h07 ;
            rom[7830] = 8'h1b ;
            rom[7831] = 8'h13 ;
            rom[7832] = 8'h00 ;
            rom[7833] = 8'hd7 ;
            rom[7834] = 8'h04 ;
            rom[7835] = 8'h04 ;
            rom[7836] = 8'hfc ;
            rom[7837] = 8'h0b ;
            rom[7838] = 8'h02 ;
            rom[7839] = 8'h01 ;
            rom[7840] = 8'h10 ;
            rom[7841] = 8'hf2 ;
            rom[7842] = 8'hd7 ;
            rom[7843] = 8'he2 ;
            rom[7844] = 8'hfd ;
            rom[7845] = 8'hf7 ;
            rom[7846] = 8'hf8 ;
            rom[7847] = 8'heb ;
            rom[7848] = 8'hfa ;
            rom[7849] = 8'hd1 ;
            rom[7850] = 8'h02 ;
            rom[7851] = 8'h08 ;
            rom[7852] = 8'h00 ;
            rom[7853] = 8'hf7 ;
            rom[7854] = 8'hf1 ;
            rom[7855] = 8'h03 ;
            rom[7856] = 8'hf7 ;
            rom[7857] = 8'h07 ;
            rom[7858] = 8'hfd ;
            rom[7859] = 8'h0b ;
            rom[7860] = 8'h03 ;
            rom[7861] = 8'h04 ;
            rom[7862] = 8'h19 ;
            rom[7863] = 8'h11 ;
            rom[7864] = 8'hf7 ;
            rom[7865] = 8'h14 ;
            rom[7866] = 8'h12 ;
            rom[7867] = 8'hfe ;
            rom[7868] = 8'h00 ;
            rom[7869] = 8'h08 ;
            rom[7870] = 8'h04 ;
            rom[7871] = 8'h02 ;
            rom[7872] = 8'h09 ;
            rom[7873] = 8'h0f ;
            rom[7874] = 8'he8 ;
            rom[7875] = 8'h0d ;
            rom[7876] = 8'h04 ;
            rom[7877] = 8'hbc ;
            rom[7878] = 8'hfb ;
            rom[7879] = 8'h09 ;
            rom[7880] = 8'h1f ;
            rom[7881] = 8'hb4 ;
            rom[7882] = 8'hdf ;
            rom[7883] = 8'h01 ;
            rom[7884] = 8'hfe ;
            rom[7885] = 8'hf4 ;
            rom[7886] = 8'he8 ;
            rom[7887] = 8'hf3 ;
            rom[7888] = 8'h26 ;
            rom[7889] = 8'hf7 ;
            rom[7890] = 8'h04 ;
            rom[7891] = 8'h05 ;
            rom[7892] = 8'hfd ;
            rom[7893] = 8'hf2 ;
            rom[7894] = 8'he8 ;
            rom[7895] = 8'h0b ;
            rom[7896] = 8'hf1 ;
            rom[7897] = 8'h09 ;
            rom[7898] = 8'hfb ;
            rom[7899] = 8'hf5 ;
            rom[7900] = 8'hd2 ;
            rom[7901] = 8'h0a ;
            rom[7902] = 8'h13 ;
            rom[7903] = 8'h0f ;
            rom[7904] = 8'hf4 ;
            rom[7905] = 8'h0c ;
            rom[7906] = 8'hc8 ;
            rom[7907] = 8'hd9 ;
            rom[7908] = 8'hfa ;
            rom[7909] = 8'hec ;
            rom[7910] = 8'hf1 ;
            rom[7911] = 8'hfe ;
            rom[7912] = 8'h1d ;
            rom[7913] = 8'he9 ;
            rom[7914] = 8'h06 ;
            rom[7915] = 8'hd8 ;
            rom[7916] = 8'he6 ;
            rom[7917] = 8'h0e ;
            rom[7918] = 8'h07 ;
            rom[7919] = 8'h05 ;
            rom[7920] = 8'h10 ;
            rom[7921] = 8'hf3 ;
            rom[7922] = 8'he5 ;
            rom[7923] = 8'h03 ;
            rom[7924] = 8'hf0 ;
            rom[7925] = 8'h14 ;
            rom[7926] = 8'hd8 ;
            rom[7927] = 8'h19 ;
            rom[7928] = 8'hcc ;
            rom[7929] = 8'hf6 ;
            rom[7930] = 8'h00 ;
            rom[7931] = 8'h12 ;
            rom[7932] = 8'h05 ;
            rom[7933] = 8'h00 ;
            rom[7934] = 8'hfe ;
            rom[7935] = 8'hf7 ;
            rom[7936] = 8'hf1 ;
            rom[7937] = 8'h15 ;
            rom[7938] = 8'hc6 ;
            rom[7939] = 8'hf8 ;
            rom[7940] = 8'h01 ;
            rom[7941] = 8'hf6 ;
            rom[7942] = 8'h12 ;
            rom[7943] = 8'h07 ;
            rom[7944] = 8'hfe ;
            rom[7945] = 8'hcd ;
            rom[7946] = 8'he5 ;
            rom[7947] = 8'h0d ;
            rom[7948] = 8'hf9 ;
            rom[7949] = 8'h1b ;
            rom[7950] = 8'hf0 ;
            rom[7951] = 8'hee ;
            rom[7952] = 8'h0a ;
            rom[7953] = 8'h26 ;
            rom[7954] = 8'h09 ;
            rom[7955] = 8'hfc ;
            rom[7956] = 8'h05 ;
            rom[7957] = 8'h10 ;
            rom[7958] = 8'hde ;
            rom[7959] = 8'h22 ;
            rom[7960] = 8'hf3 ;
            rom[7961] = 8'hea ;
            rom[7962] = 8'h08 ;
            rom[7963] = 8'h00 ;
            rom[7964] = 8'hf3 ;
            rom[7965] = 8'hd5 ;
            rom[7966] = 8'h08 ;
            rom[7967] = 8'h1c ;
            rom[7968] = 8'hbe ;
            rom[7969] = 8'hf5 ;
            rom[7970] = 8'he9 ;
            rom[7971] = 8'h10 ;
            rom[7972] = 8'h09 ;
            rom[7973] = 8'hf0 ;
            rom[7974] = 8'hf8 ;
            rom[7975] = 8'h17 ;
            rom[7976] = 8'he6 ;
            rom[7977] = 8'he5 ;
            rom[7978] = 8'he9 ;
            rom[7979] = 8'hea ;
            rom[7980] = 8'hf6 ;
            rom[7981] = 8'h08 ;
            rom[7982] = 8'he9 ;
            rom[7983] = 8'hf1 ;
            rom[7984] = 8'h0a ;
            rom[7985] = 8'h2a ;
            rom[7986] = 8'hef ;
            rom[7987] = 8'hfa ;
            rom[7988] = 8'hfc ;
            rom[7989] = 8'hf5 ;
            rom[7990] = 8'h23 ;
            rom[7991] = 8'h1f ;
            rom[7992] = 8'hd0 ;
            rom[7993] = 8'hf0 ;
            rom[7994] = 8'hfd ;
            rom[7995] = 8'h1e ;
            rom[7996] = 8'he5 ;
            rom[7997] = 8'hf1 ;
            rom[7998] = 8'hfc ;
            rom[7999] = 8'hf8 ;
            rom[8000] = 8'h25 ;
            rom[8001] = 8'h08 ;
            rom[8002] = 8'h0c ;
            rom[8003] = 8'hf1 ;
            rom[8004] = 8'h13 ;
            rom[8005] = 8'h1d ;
            rom[8006] = 8'h06 ;
            rom[8007] = 8'hd8 ;
            rom[8008] = 8'hfc ;
            rom[8009] = 8'h04 ;
            rom[8010] = 8'hf3 ;
            rom[8011] = 8'h06 ;
            rom[8012] = 8'hee ;
            rom[8013] = 8'he0 ;
            rom[8014] = 8'h03 ;
            rom[8015] = 8'hdc ;
            rom[8016] = 8'hf5 ;
            rom[8017] = 8'h38 ;
            rom[8018] = 8'hfd ;
            rom[8019] = 8'hea ;
            rom[8020] = 8'hbe ;
            rom[8021] = 8'hd9 ;
            rom[8022] = 8'h11 ;
            rom[8023] = 8'h01 ;
            rom[8024] = 8'hf3 ;
            rom[8025] = 8'hf5 ;
            rom[8026] = 8'h0b ;
            rom[8027] = 8'he9 ;
            rom[8028] = 8'h0c ;
            rom[8029] = 8'h1d ;
            rom[8030] = 8'h15 ;
            rom[8031] = 8'h1c ;
            rom[8032] = 8'hf4 ;
            rom[8033] = 8'h05 ;
            rom[8034] = 8'h0f ;
            rom[8035] = 8'h00 ;
            rom[8036] = 8'h0f ;
            rom[8037] = 8'h12 ;
            rom[8038] = 8'h28 ;
            rom[8039] = 8'heb ;
            rom[8040] = 8'h03 ;
            rom[8041] = 8'hdf ;
            rom[8042] = 8'h24 ;
            rom[8043] = 8'h0b ;
            rom[8044] = 8'hd0 ;
            rom[8045] = 8'h02 ;
            rom[8046] = 8'h03 ;
            rom[8047] = 8'hee ;
            rom[8048] = 8'h1b ;
            rom[8049] = 8'hfa ;
            rom[8050] = 8'hed ;
            rom[8051] = 8'he5 ;
            rom[8052] = 8'hee ;
            rom[8053] = 8'h05 ;
            rom[8054] = 8'he3 ;
            rom[8055] = 8'h21 ;
            rom[8056] = 8'hfb ;
            rom[8057] = 8'h07 ;
            rom[8058] = 8'hfd ;
            rom[8059] = 8'hf4 ;
            rom[8060] = 8'h05 ;
            rom[8061] = 8'hf6 ;
            rom[8062] = 8'he5 ;
            rom[8063] = 8'h15 ;
            rom[8064] = 8'hfb ;
            rom[8065] = 8'h09 ;
            rom[8066] = 8'he7 ;
            rom[8067] = 8'hf2 ;
            rom[8068] = 8'h21 ;
            rom[8069] = 8'h09 ;
            rom[8070] = 8'he5 ;
            rom[8071] = 8'hd8 ;
            rom[8072] = 8'hf6 ;
            rom[8073] = 8'h0f ;
            rom[8074] = 8'h03 ;
            rom[8075] = 8'h18 ;
            rom[8076] = 8'h14 ;
            rom[8077] = 8'hf0 ;
            rom[8078] = 8'h06 ;
            rom[8079] = 8'hfe ;
            rom[8080] = 8'h03 ;
            rom[8081] = 8'h13 ;
            rom[8082] = 8'hfe ;
            rom[8083] = 8'h15 ;
            rom[8084] = 8'h0b ;
            rom[8085] = 8'hf0 ;
            rom[8086] = 8'h0c ;
            rom[8087] = 8'h09 ;
            rom[8088] = 8'he0 ;
            rom[8089] = 8'hf5 ;
            rom[8090] = 8'hf6 ;
            rom[8091] = 8'h1e ;
            rom[8092] = 8'h0c ;
            rom[8093] = 8'hfd ;
            rom[8094] = 8'hef ;
            rom[8095] = 8'hf9 ;
            rom[8096] = 8'hda ;
            rom[8097] = 8'hfe ;
            rom[8098] = 8'hf4 ;
            rom[8099] = 8'hf7 ;
            rom[8100] = 8'h16 ;
            rom[8101] = 8'hf3 ;
            rom[8102] = 8'h04 ;
            rom[8103] = 8'h1c ;
            rom[8104] = 8'h03 ;
            rom[8105] = 8'he4 ;
            rom[8106] = 8'hf2 ;
            rom[8107] = 8'h05 ;
            rom[8108] = 8'h13 ;
            rom[8109] = 8'h32 ;
            rom[8110] = 8'h11 ;
            rom[8111] = 8'he5 ;
            rom[8112] = 8'h18 ;
            rom[8113] = 8'he5 ;
            rom[8114] = 8'hf2 ;
            rom[8115] = 8'hf5 ;
            rom[8116] = 8'h26 ;
            rom[8117] = 8'hf4 ;
            rom[8118] = 8'h09 ;
            rom[8119] = 8'h0c ;
            rom[8120] = 8'hfc ;
            rom[8121] = 8'h04 ;
            rom[8122] = 8'h07 ;
            rom[8123] = 8'he6 ;
            rom[8124] = 8'hf7 ;
            rom[8125] = 8'hd9 ;
            rom[8126] = 8'h10 ;
            rom[8127] = 8'hed ;
            rom[8128] = 8'h1b ;
            rom[8129] = 8'hff ;
            rom[8130] = 8'hf1 ;
            rom[8131] = 8'hfe ;
            rom[8132] = 8'h21 ;
            rom[8133] = 8'hff ;
            rom[8134] = 8'h00 ;
            rom[8135] = 8'h1f ;
            rom[8136] = 8'h14 ;
            rom[8137] = 8'he5 ;
            rom[8138] = 8'h05 ;
            rom[8139] = 8'hfd ;
            rom[8140] = 8'hfb ;
            rom[8141] = 8'he7 ;
            rom[8142] = 8'h15 ;
            rom[8143] = 8'he0 ;
            rom[8144] = 8'hf3 ;
            rom[8145] = 8'h22 ;
            rom[8146] = 8'hf0 ;
            rom[8147] = 8'hd8 ;
            rom[8148] = 8'hef ;
            rom[8149] = 8'h02 ;
            rom[8150] = 8'h12 ;
            rom[8151] = 8'hfc ;
            rom[8152] = 8'hea ;
            rom[8153] = 8'h12 ;
            rom[8154] = 8'h0c ;
            rom[8155] = 8'h0a ;
            rom[8156] = 8'h0a ;
            rom[8157] = 8'hf4 ;
            rom[8158] = 8'he2 ;
            rom[8159] = 8'h1f ;
            rom[8160] = 8'h06 ;
            rom[8161] = 8'h08 ;
            rom[8162] = 8'h03 ;
            rom[8163] = 8'h0d ;
            rom[8164] = 8'h0d ;
            rom[8165] = 8'hf2 ;
            rom[8166] = 8'h0b ;
            rom[8167] = 8'hd0 ;
            rom[8168] = 8'hf1 ;
            rom[8169] = 8'h0b ;
            rom[8170] = 8'h17 ;
            rom[8171] = 8'h0c ;
            rom[8172] = 8'hf3 ;
            rom[8173] = 8'h15 ;
            rom[8174] = 8'h06 ;
            rom[8175] = 8'h10 ;
            rom[8176] = 8'h00 ;
            rom[8177] = 8'hf3 ;
            rom[8178] = 8'hec ;
            rom[8179] = 8'hf2 ;
            rom[8180] = 8'he6 ;
            rom[8181] = 8'h08 ;
            rom[8182] = 8'h10 ;
            rom[8183] = 8'hfb ;
            rom[8184] = 8'hd4 ;
            rom[8185] = 8'h09 ;
            rom[8186] = 8'h2e ;
            rom[8187] = 8'hf7 ;
            rom[8188] = 8'h04 ;
            rom[8189] = 8'h10 ;
            rom[8190] = 8'h06 ;
            rom[8191] = 8'h26 ;
            rom[8192] = 8'h18 ;
            rom[8193] = 8'h0c ;
            rom[8194] = 8'he8 ;
            rom[8195] = 8'h05 ;
            rom[8196] = 8'hf4 ;
            rom[8197] = 8'hfd ;
            rom[8198] = 8'hf4 ;
            rom[8199] = 8'hc4 ;
            rom[8200] = 8'hfc ;
            rom[8201] = 8'hfc ;
            rom[8202] = 8'hfa ;
            rom[8203] = 8'hef ;
            rom[8204] = 8'ha4 ;
            rom[8205] = 8'he0 ;
            rom[8206] = 8'h1c ;
            rom[8207] = 8'hdd ;
            rom[8208] = 8'hff ;
            rom[8209] = 8'hf4 ;
            rom[8210] = 8'hfa ;
            rom[8211] = 8'hfd ;
            rom[8212] = 8'hde ;
            rom[8213] = 8'h0c ;
            rom[8214] = 8'hf7 ;
            rom[8215] = 8'h05 ;
            rom[8216] = 8'he8 ;
            rom[8217] = 8'h04 ;
            rom[8218] = 8'h0a ;
            rom[8219] = 8'hec ;
            rom[8220] = 8'h01 ;
            rom[8221] = 8'h09 ;
            rom[8222] = 8'hf1 ;
            rom[8223] = 8'h17 ;
            rom[8224] = 8'h13 ;
            rom[8225] = 8'h03 ;
            rom[8226] = 8'hf9 ;
            rom[8227] = 8'hf7 ;
            rom[8228] = 8'hea ;
            rom[8229] = 8'h21 ;
            rom[8230] = 8'hec ;
            rom[8231] = 8'hde ;
            rom[8232] = 8'hf9 ;
            rom[8233] = 8'hed ;
            rom[8234] = 8'hee ;
            rom[8235] = 8'h09 ;
            rom[8236] = 8'h16 ;
            rom[8237] = 8'hf1 ;
            rom[8238] = 8'h13 ;
            rom[8239] = 8'he1 ;
            rom[8240] = 8'he4 ;
            rom[8241] = 8'h0a ;
            rom[8242] = 8'h1e ;
            rom[8243] = 8'hd9 ;
            rom[8244] = 8'hf3 ;
            rom[8245] = 8'hf1 ;
            rom[8246] = 8'he4 ;
            rom[8247] = 8'hd9 ;
            rom[8248] = 8'hee ;
            rom[8249] = 8'h10 ;
            rom[8250] = 8'hed ;
            rom[8251] = 8'hda ;
            rom[8252] = 8'hfd ;
            rom[8253] = 8'h01 ;
            rom[8254] = 8'hf3 ;
            rom[8255] = 8'he2 ;
            rom[8256] = 8'h0a ;
            rom[8257] = 8'he7 ;
            rom[8258] = 8'h09 ;
            rom[8259] = 8'hd1 ;
            rom[8260] = 8'h11 ;
            rom[8261] = 8'h1c ;
            rom[8262] = 8'hf1 ;
            rom[8263] = 8'hee ;
            rom[8264] = 8'he4 ;
            rom[8265] = 8'h15 ;
            rom[8266] = 8'h05 ;
            rom[8267] = 8'hc3 ;
            rom[8268] = 8'h10 ;
            rom[8269] = 8'hec ;
            rom[8270] = 8'hd6 ;
            rom[8271] = 8'hed ;
            rom[8272] = 8'h12 ;
            rom[8273] = 8'hfa ;
            rom[8274] = 8'h1a ;
            rom[8275] = 8'h04 ;
            rom[8276] = 8'he7 ;
            rom[8277] = 8'he5 ;
            rom[8278] = 8'hfb ;
            rom[8279] = 8'h17 ;
            rom[8280] = 8'hef ;
            rom[8281] = 8'heb ;
            rom[8282] = 8'hcf ;
            rom[8283] = 8'hd8 ;
            rom[8284] = 8'hfa ;
            rom[8285] = 8'h16 ;
            rom[8286] = 8'h08 ;
            rom[8287] = 8'hf1 ;
            rom[8288] = 8'hfe ;
            rom[8289] = 8'hea ;
            rom[8290] = 8'hf2 ;
            rom[8291] = 8'he2 ;
            rom[8292] = 8'hff ;
            rom[8293] = 8'h17 ;
            rom[8294] = 8'hfa ;
            rom[8295] = 8'he8 ;
            rom[8296] = 8'h10 ;
            rom[8297] = 8'he8 ;
            rom[8298] = 8'h0a ;
            rom[8299] = 8'hfd ;
            rom[8300] = 8'hf9 ;
            rom[8301] = 8'hf8 ;
            rom[8302] = 8'hdf ;
            rom[8303] = 8'hfc ;
            rom[8304] = 8'he4 ;
            rom[8305] = 8'hd8 ;
            rom[8306] = 8'h1d ;
            rom[8307] = 8'hfd ;
            rom[8308] = 8'hbd ;
            rom[8309] = 8'h01 ;
            rom[8310] = 8'h0b ;
            rom[8311] = 8'hfe ;
            rom[8312] = 8'h19 ;
            rom[8313] = 8'he7 ;
            rom[8314] = 8'hdf ;
            rom[8315] = 8'h21 ;
            rom[8316] = 8'hfd ;
            rom[8317] = 8'he4 ;
            rom[8318] = 8'h17 ;
            rom[8319] = 8'h06 ;
            rom[8320] = 8'h0b ;
            rom[8321] = 8'hef ;
            rom[8322] = 8'h13 ;
            rom[8323] = 8'h19 ;
            rom[8324] = 8'h08 ;
            rom[8325] = 8'hc4 ;
            rom[8326] = 8'hd6 ;
            rom[8327] = 8'h1a ;
            rom[8328] = 8'h1b ;
            rom[8329] = 8'hdb ;
            rom[8330] = 8'h0a ;
            rom[8331] = 8'h0e ;
            rom[8332] = 8'h03 ;
            rom[8333] = 8'hda ;
            rom[8334] = 8'hff ;
            rom[8335] = 8'hfc ;
            rom[8336] = 8'hfe ;
            rom[8337] = 8'h16 ;
            rom[8338] = 8'he5 ;
            rom[8339] = 8'he5 ;
            rom[8340] = 8'h05 ;
            rom[8341] = 8'h0b ;
            rom[8342] = 8'h03 ;
            rom[8343] = 8'hea ;
            rom[8344] = 8'hee ;
            rom[8345] = 8'h10 ;
            rom[8346] = 8'hc8 ;
            rom[8347] = 8'h21 ;
            rom[8348] = 8'hec ;
            rom[8349] = 8'hfe ;
            rom[8350] = 8'h0a ;
            rom[8351] = 8'hfa ;
            rom[8352] = 8'h00 ;
            rom[8353] = 8'hd3 ;
            rom[8354] = 8'hfa ;
            rom[8355] = 8'h02 ;
            rom[8356] = 8'hf8 ;
            rom[8357] = 8'h01 ;
            rom[8358] = 8'hf8 ;
            rom[8359] = 8'hdb ;
            rom[8360] = 8'hea ;
            rom[8361] = 8'hfa ;
            rom[8362] = 8'h03 ;
            rom[8363] = 8'h12 ;
            rom[8364] = 8'hf4 ;
            rom[8365] = 8'he7 ;
            rom[8366] = 8'he4 ;
            rom[8367] = 8'hfd ;
            rom[8368] = 8'h05 ;
            rom[8369] = 8'hfc ;
            rom[8370] = 8'hfa ;
            rom[8371] = 8'hf9 ;
            rom[8372] = 8'hfa ;
            rom[8373] = 8'hfe ;
            rom[8374] = 8'h0a ;
            rom[8375] = 8'hf3 ;
            rom[8376] = 8'he6 ;
            rom[8377] = 8'he0 ;
            rom[8378] = 8'h17 ;
            rom[8379] = 8'he1 ;
            rom[8380] = 8'hf2 ;
            rom[8381] = 8'he9 ;
            rom[8382] = 8'h3a ;
            rom[8383] = 8'hd1 ;
            rom[8384] = 8'h1b ;
            rom[8385] = 8'h07 ;
            rom[8386] = 8'hf5 ;
            rom[8387] = 8'h15 ;
            rom[8388] = 8'h07 ;
            rom[8389] = 8'hc7 ;
            rom[8390] = 8'hdf ;
            rom[8391] = 8'hf7 ;
            rom[8392] = 8'h16 ;
            rom[8393] = 8'he4 ;
            rom[8394] = 8'h08 ;
            rom[8395] = 8'hf6 ;
            rom[8396] = 8'hdb ;
            rom[8397] = 8'he7 ;
            rom[8398] = 8'h22 ;
            rom[8399] = 8'h06 ;
            rom[8400] = 8'hf2 ;
            rom[8401] = 8'h0f ;
            rom[8402] = 8'hfe ;
            rom[8403] = 8'he0 ;
            rom[8404] = 8'h1c ;
            rom[8405] = 8'he0 ;
            rom[8406] = 8'hdf ;
            rom[8407] = 8'hcb ;
            rom[8408] = 8'h06 ;
            rom[8409] = 8'h16 ;
            rom[8410] = 8'hfc ;
            rom[8411] = 8'h09 ;
            rom[8412] = 8'h14 ;
            rom[8413] = 8'h11 ;
            rom[8414] = 8'h08 ;
            rom[8415] = 8'hf7 ;
            rom[8416] = 8'h19 ;
            rom[8417] = 8'h06 ;
            rom[8418] = 8'h0d ;
            rom[8419] = 8'hfd ;
            rom[8420] = 8'hf7 ;
            rom[8421] = 8'h02 ;
            rom[8422] = 8'h12 ;
            rom[8423] = 8'hef ;
            rom[8424] = 8'he2 ;
            rom[8425] = 8'hf7 ;
            rom[8426] = 8'hd6 ;
            rom[8427] = 8'h09 ;
            rom[8428] = 8'h10 ;
            rom[8429] = 8'hda ;
            rom[8430] = 8'hf9 ;
            rom[8431] = 8'hdd ;
            rom[8432] = 8'hf7 ;
            rom[8433] = 8'he4 ;
            rom[8434] = 8'h0c ;
            rom[8435] = 8'hda ;
            rom[8436] = 8'h0e ;
            rom[8437] = 8'he3 ;
            rom[8438] = 8'hfb ;
            rom[8439] = 8'he7 ;
            rom[8440] = 8'h00 ;
            rom[8441] = 8'h10 ;
            rom[8442] = 8'h17 ;
            rom[8443] = 8'h03 ;
            rom[8444] = 8'he5 ;
            rom[8445] = 8'hea ;
            rom[8446] = 8'h06 ;
            rom[8447] = 8'hd2 ;
            rom[8448] = 8'h29 ;
            rom[8449] = 8'hf5 ;
            rom[8450] = 8'hf4 ;
            rom[8451] = 8'he9 ;
            rom[8452] = 8'h14 ;
            rom[8453] = 8'hf3 ;
            rom[8454] = 8'h0e ;
            rom[8455] = 8'h12 ;
            rom[8456] = 8'hf2 ;
            rom[8457] = 8'hf1 ;
            rom[8458] = 8'hf9 ;
            rom[8459] = 8'hde ;
            rom[8460] = 8'hda ;
            rom[8461] = 8'hed ;
            rom[8462] = 8'h09 ;
            rom[8463] = 8'h0c ;
            rom[8464] = 8'h14 ;
            rom[8465] = 8'heb ;
            rom[8466] = 8'h14 ;
            rom[8467] = 8'h11 ;
            rom[8468] = 8'he3 ;
            rom[8469] = 8'hf7 ;
            rom[8470] = 8'hef ;
            rom[8471] = 8'h16 ;
            rom[8472] = 8'h04 ;
            rom[8473] = 8'h03 ;
            rom[8474] = 8'hf3 ;
            rom[8475] = 8'hff ;
            rom[8476] = 8'h04 ;
            rom[8477] = 8'h01 ;
            rom[8478] = 8'h04 ;
            rom[8479] = 8'h01 ;
            rom[8480] = 8'hfc ;
            rom[8481] = 8'hef ;
            rom[8482] = 8'he5 ;
            rom[8483] = 8'hef ;
            rom[8484] = 8'h1b ;
            rom[8485] = 8'h1b ;
            rom[8486] = 8'hd1 ;
            rom[8487] = 8'hfb ;
            rom[8488] = 8'h0b ;
            rom[8489] = 8'hf3 ;
            rom[8490] = 8'hde ;
            rom[8491] = 8'hf1 ;
            rom[8492] = 8'hcc ;
            rom[8493] = 8'h01 ;
            rom[8494] = 8'hca ;
            rom[8495] = 8'h0b ;
            rom[8496] = 8'hf1 ;
            rom[8497] = 8'h20 ;
            rom[8498] = 8'h02 ;
            rom[8499] = 8'hd7 ;
            rom[8500] = 8'h03 ;
            rom[8501] = 8'hec ;
            rom[8502] = 8'hd7 ;
            rom[8503] = 8'hed ;
            rom[8504] = 8'h1a ;
            rom[8505] = 8'hfa ;
            rom[8506] = 8'hef ;
            rom[8507] = 8'h0b ;
            rom[8508] = 8'h00 ;
            rom[8509] = 8'hf4 ;
            rom[8510] = 8'hea ;
            rom[8511] = 8'h04 ;
            rom[8512] = 8'h3e ;
            rom[8513] = 8'heb ;
            rom[8514] = 8'hfd ;
            rom[8515] = 8'h0e ;
            rom[8516] = 8'hc3 ;
            rom[8517] = 8'he5 ;
            rom[8518] = 8'hf4 ;
            rom[8519] = 8'h04 ;
            rom[8520] = 8'h08 ;
            rom[8521] = 8'hce ;
            rom[8522] = 8'h12 ;
            rom[8523] = 8'h23 ;
            rom[8524] = 8'h0c ;
            rom[8525] = 8'hf0 ;
            rom[8526] = 8'he8 ;
            rom[8527] = 8'hf0 ;
            rom[8528] = 8'hff ;
            rom[8529] = 8'h0b ;
            rom[8530] = 8'h00 ;
            rom[8531] = 8'he6 ;
            rom[8532] = 8'hf9 ;
            rom[8533] = 8'hfd ;
            rom[8534] = 8'h26 ;
            rom[8535] = 8'h06 ;
            rom[8536] = 8'h11 ;
            rom[8537] = 8'hf4 ;
            rom[8538] = 8'hf3 ;
            rom[8539] = 8'he2 ;
            rom[8540] = 8'h01 ;
            rom[8541] = 8'hf0 ;
            rom[8542] = 8'h1f ;
            rom[8543] = 8'h19 ;
            rom[8544] = 8'h08 ;
            rom[8545] = 8'h15 ;
            rom[8546] = 8'hcb ;
            rom[8547] = 8'hdb ;
            rom[8548] = 8'hf1 ;
            rom[8549] = 8'h1b ;
            rom[8550] = 8'h06 ;
            rom[8551] = 8'h26 ;
            rom[8552] = 8'hcc ;
            rom[8553] = 8'hfe ;
            rom[8554] = 8'h15 ;
            rom[8555] = 8'hd4 ;
            rom[8556] = 8'he5 ;
            rom[8557] = 8'heb ;
            rom[8558] = 8'h21 ;
            rom[8559] = 8'hef ;
            rom[8560] = 8'h0f ;
            rom[8561] = 8'hd6 ;
            rom[8562] = 8'hd7 ;
            rom[8563] = 8'hfd ;
            rom[8564] = 8'hdf ;
            rom[8565] = 8'hf1 ;
            rom[8566] = 8'hf4 ;
            rom[8567] = 8'hef ;
            rom[8568] = 8'hfc ;
            rom[8569] = 8'h07 ;
            rom[8570] = 8'h0d ;
            rom[8571] = 8'h16 ;
            rom[8572] = 8'h14 ;
            rom[8573] = 8'h07 ;
            rom[8574] = 8'h07 ;
            rom[8575] = 8'h1f ;
            rom[8576] = 8'hfc ;
            rom[8577] = 8'hfc ;
            rom[8578] = 8'h01 ;
            rom[8579] = 8'h09 ;
            rom[8580] = 8'h0e ;
            rom[8581] = 8'hf2 ;
            rom[8582] = 8'h0a ;
            rom[8583] = 8'hfa ;
            rom[8584] = 8'h0f ;
            rom[8585] = 8'hee ;
            rom[8586] = 8'h1f ;
            rom[8587] = 8'hfc ;
            rom[8588] = 8'hf6 ;
            rom[8589] = 8'h0a ;
            rom[8590] = 8'h02 ;
            rom[8591] = 8'h13 ;
            rom[8592] = 8'h12 ;
            rom[8593] = 8'h1a ;
            rom[8594] = 8'hf6 ;
            rom[8595] = 8'h18 ;
            rom[8596] = 8'h04 ;
            rom[8597] = 8'h06 ;
            rom[8598] = 8'h06 ;
            rom[8599] = 8'hda ;
            rom[8600] = 8'hb8 ;
            rom[8601] = 8'hf9 ;
            rom[8602] = 8'he8 ;
            rom[8603] = 8'h13 ;
            rom[8604] = 8'ha6 ;
            rom[8605] = 8'h01 ;
            rom[8606] = 8'h03 ;
            rom[8607] = 8'h05 ;
            rom[8608] = 8'h0c ;
            rom[8609] = 8'he5 ;
            rom[8610] = 8'hff ;
            rom[8611] = 8'hec ;
            rom[8612] = 8'hf1 ;
            rom[8613] = 8'h21 ;
            rom[8614] = 8'he7 ;
            rom[8615] = 8'h14 ;
            rom[8616] = 8'h02 ;
            rom[8617] = 8'h0e ;
            rom[8618] = 8'h05 ;
            rom[8619] = 8'h0d ;
            rom[8620] = 8'h1a ;
            rom[8621] = 8'hbc ;
            rom[8622] = 8'hfb ;
            rom[8623] = 8'h03 ;
            rom[8624] = 8'hfb ;
            rom[8625] = 8'h05 ;
            rom[8626] = 8'hc5 ;
            rom[8627] = 8'h1c ;
            rom[8628] = 8'h14 ;
            rom[8629] = 8'he3 ;
            rom[8630] = 8'hf8 ;
            rom[8631] = 8'hf2 ;
            rom[8632] = 8'hd9 ;
            rom[8633] = 8'h15 ;
            rom[8634] = 8'he3 ;
            rom[8635] = 8'h1f ;
            rom[8636] = 8'hd6 ;
            rom[8637] = 8'hcf ;
            rom[8638] = 8'h27 ;
            rom[8639] = 8'hc3 ;
            rom[8640] = 8'h29 ;
            rom[8641] = 8'hee ;
            rom[8642] = 8'h34 ;
            rom[8643] = 8'hde ;
            rom[8644] = 8'he7 ;
            rom[8645] = 8'h19 ;
            rom[8646] = 8'hfe ;
            rom[8647] = 8'hf3 ;
            rom[8648] = 8'hff ;
            rom[8649] = 8'hf3 ;
            rom[8650] = 8'h09 ;
            rom[8651] = 8'hd9 ;
            rom[8652] = 8'h07 ;
            rom[8653] = 8'hf5 ;
            rom[8654] = 8'h01 ;
            rom[8655] = 8'h04 ;
            rom[8656] = 8'hf8 ;
            rom[8657] = 8'h10 ;
            rom[8658] = 8'h22 ;
            rom[8659] = 8'h03 ;
            rom[8660] = 8'hfe ;
            rom[8661] = 8'h09 ;
            rom[8662] = 8'h00 ;
            rom[8663] = 8'h05 ;
            rom[8664] = 8'he7 ;
            rom[8665] = 8'h03 ;
            rom[8666] = 8'he8 ;
            rom[8667] = 8'h01 ;
            rom[8668] = 8'h0a ;
            rom[8669] = 8'h03 ;
            rom[8670] = 8'h00 ;
            rom[8671] = 8'hfd ;
            rom[8672] = 8'h21 ;
            rom[8673] = 8'hf1 ;
            rom[8674] = 8'h17 ;
            rom[8675] = 8'hfc ;
            rom[8676] = 8'h02 ;
            rom[8677] = 8'h28 ;
            rom[8678] = 8'h15 ;
            rom[8679] = 8'h03 ;
            rom[8680] = 8'hfc ;
            rom[8681] = 8'h01 ;
            rom[8682] = 8'hfd ;
            rom[8683] = 8'h08 ;
            rom[8684] = 8'h15 ;
            rom[8685] = 8'hdb ;
            rom[8686] = 8'hff ;
            rom[8687] = 8'he1 ;
            rom[8688] = 8'h01 ;
            rom[8689] = 8'he1 ;
            rom[8690] = 8'hef ;
            rom[8691] = 8'hd8 ;
            rom[8692] = 8'h16 ;
            rom[8693] = 8'h00 ;
            rom[8694] = 8'he8 ;
            rom[8695] = 8'hf0 ;
            rom[8696] = 8'h0b ;
            rom[8697] = 8'hf2 ;
            rom[8698] = 8'heb ;
            rom[8699] = 8'hfa ;
            rom[8700] = 8'hee ;
            rom[8701] = 8'hc3 ;
            rom[8702] = 8'h21 ;
            rom[8703] = 8'hfc ;
            rom[8704] = 8'h08 ;
            rom[8705] = 8'h0f ;
            rom[8706] = 8'hea ;
            rom[8707] = 8'hd2 ;
            rom[8708] = 8'hf5 ;
            rom[8709] = 8'h11 ;
            rom[8710] = 8'hf5 ;
            rom[8711] = 8'hed ;
            rom[8712] = 8'h03 ;
            rom[8713] = 8'he3 ;
            rom[8714] = 8'he3 ;
            rom[8715] = 8'hd2 ;
            rom[8716] = 8'h00 ;
            rom[8717] = 8'hec ;
            rom[8718] = 8'hfe ;
            rom[8719] = 8'h09 ;
            rom[8720] = 8'h20 ;
            rom[8721] = 8'h0a ;
            rom[8722] = 8'h01 ;
            rom[8723] = 8'hd8 ;
            rom[8724] = 8'haa ;
            rom[8725] = 8'hdc ;
            rom[8726] = 8'h08 ;
            rom[8727] = 8'h1c ;
            rom[8728] = 8'h07 ;
            rom[8729] = 8'hed ;
            rom[8730] = 8'hfd ;
            rom[8731] = 8'hd3 ;
            rom[8732] = 8'hf1 ;
            rom[8733] = 8'h0e ;
            rom[8734] = 8'hfc ;
            rom[8735] = 8'hb9 ;
            rom[8736] = 8'h12 ;
            rom[8737] = 8'hd8 ;
            rom[8738] = 8'hec ;
            rom[8739] = 8'hfc ;
            rom[8740] = 8'h06 ;
            rom[8741] = 8'h35 ;
            rom[8742] = 8'hdf ;
            rom[8743] = 8'h13 ;
            rom[8744] = 8'h0d ;
            rom[8745] = 8'hc5 ;
            rom[8746] = 8'h0d ;
            rom[8747] = 8'hc9 ;
            rom[8748] = 8'h05 ;
            rom[8749] = 8'h0a ;
            rom[8750] = 8'hf8 ;
            rom[8751] = 8'h09 ;
            rom[8752] = 8'hff ;
            rom[8753] = 8'hc3 ;
            rom[8754] = 8'h16 ;
            rom[8755] = 8'h09 ;
            rom[8756] = 8'ha7 ;
            rom[8757] = 8'hf6 ;
            rom[8758] = 8'hfc ;
            rom[8759] = 8'hfe ;
            rom[8760] = 8'h12 ;
            rom[8761] = 8'h01 ;
            rom[8762] = 8'h02 ;
            rom[8763] = 8'hfd ;
            rom[8764] = 8'hfc ;
            rom[8765] = 8'hd8 ;
            rom[8766] = 8'hfb ;
            rom[8767] = 8'hdf ;
            rom[8768] = 8'h13 ;
            rom[8769] = 8'h09 ;
            rom[8770] = 8'h22 ;
            rom[8771] = 8'hcc ;
            rom[8772] = 8'h14 ;
            rom[8773] = 8'h14 ;
            rom[8774] = 8'hf7 ;
            rom[8775] = 8'he6 ;
            rom[8776] = 8'hfb ;
            rom[8777] = 8'hef ;
            rom[8778] = 8'h14 ;
            rom[8779] = 8'hc8 ;
            rom[8780] = 8'h02 ;
            rom[8781] = 8'he1 ;
            rom[8782] = 8'he4 ;
            rom[8783] = 8'hd8 ;
            rom[8784] = 8'h0c ;
            rom[8785] = 8'h11 ;
            rom[8786] = 8'hf9 ;
            rom[8787] = 8'hed ;
            rom[8788] = 8'he6 ;
            rom[8789] = 8'hf2 ;
            rom[8790] = 8'he1 ;
            rom[8791] = 8'h28 ;
            rom[8792] = 8'hf1 ;
            rom[8793] = 8'he5 ;
            rom[8794] = 8'hd9 ;
            rom[8795] = 8'hd8 ;
            rom[8796] = 8'h11 ;
            rom[8797] = 8'h0e ;
            rom[8798] = 8'h09 ;
            rom[8799] = 8'hc4 ;
            rom[8800] = 8'hfa ;
            rom[8801] = 8'hec ;
            rom[8802] = 8'h18 ;
            rom[8803] = 8'he8 ;
            rom[8804] = 8'h11 ;
            rom[8805] = 8'h34 ;
            rom[8806] = 8'he5 ;
            rom[8807] = 8'hec ;
            rom[8808] = 8'h0a ;
            rom[8809] = 8'hd4 ;
            rom[8810] = 8'h1f ;
            rom[8811] = 8'h03 ;
            rom[8812] = 8'h00 ;
            rom[8813] = 8'he0 ;
            rom[8814] = 8'hd1 ;
            rom[8815] = 8'h06 ;
            rom[8816] = 8'hdc ;
            rom[8817] = 8'hda ;
            rom[8818] = 8'h14 ;
            rom[8819] = 8'h1a ;
            rom[8820] = 8'hbb ;
            rom[8821] = 8'hed ;
            rom[8822] = 8'h0e ;
            rom[8823] = 8'hea ;
            rom[8824] = 8'h2a ;
            rom[8825] = 8'hf8 ;
            rom[8826] = 8'he4 ;
            rom[8827] = 8'h0e ;
            rom[8828] = 8'hf9 ;
            rom[8829] = 8'he2 ;
            rom[8830] = 8'h03 ;
            rom[8831] = 8'h07 ;
            rom[8832] = 8'h0b ;
            rom[8833] = 8'hcf ;
            rom[8834] = 8'h06 ;
            rom[8835] = 8'h02 ;
            rom[8836] = 8'h02 ;
            rom[8837] = 8'h05 ;
            rom[8838] = 8'h13 ;
            rom[8839] = 8'hcf ;
            rom[8840] = 8'hfe ;
            rom[8841] = 8'hf8 ;
            rom[8842] = 8'h12 ;
            rom[8843] = 8'h1c ;
            rom[8844] = 8'hfb ;
            rom[8845] = 8'hff ;
            rom[8846] = 8'hf9 ;
            rom[8847] = 8'hfe ;
            rom[8848] = 8'hf5 ;
            rom[8849] = 8'h15 ;
            rom[8850] = 8'h07 ;
            rom[8851] = 8'hf7 ;
            rom[8852] = 8'hff ;
            rom[8853] = 8'h0b ;
            rom[8854] = 8'heb ;
            rom[8855] = 8'hf1 ;
            rom[8856] = 8'h1b ;
            rom[8857] = 8'hfc ;
            rom[8858] = 8'hf0 ;
            rom[8859] = 8'ha6 ;
            rom[8860] = 8'h04 ;
            rom[8861] = 8'h04 ;
            rom[8862] = 8'h13 ;
            rom[8863] = 8'hfa ;
            rom[8864] = 8'h00 ;
            rom[8865] = 8'h00 ;
            rom[8866] = 8'h00 ;
            rom[8867] = 8'hfd ;
            rom[8868] = 8'hf7 ;
            rom[8869] = 8'h17 ;
            rom[8870] = 8'h0a ;
            rom[8871] = 8'h06 ;
            rom[8872] = 8'hc5 ;
            rom[8873] = 8'h05 ;
            rom[8874] = 8'h03 ;
            rom[8875] = 8'he4 ;
            rom[8876] = 8'h49 ;
            rom[8877] = 8'h05 ;
            rom[8878] = 8'h1c ;
            rom[8879] = 8'h20 ;
            rom[8880] = 8'hce ;
            rom[8881] = 8'hfc ;
            rom[8882] = 8'h0d ;
            rom[8883] = 8'hfe ;
            rom[8884] = 8'hfb ;
            rom[8885] = 8'h00 ;
            rom[8886] = 8'h08 ;
            rom[8887] = 8'hd6 ;
            rom[8888] = 8'h02 ;
            rom[8889] = 8'hfc ;
            rom[8890] = 8'hef ;
            rom[8891] = 8'h26 ;
            rom[8892] = 8'h1a ;
            rom[8893] = 8'hfe ;
            rom[8894] = 8'h11 ;
            rom[8895] = 8'h1a ;
            rom[8896] = 8'h05 ;
            rom[8897] = 8'h14 ;
            rom[8898] = 8'h06 ;
            rom[8899] = 8'hf5 ;
            rom[8900] = 8'h13 ;
            rom[8901] = 8'hfd ;
            rom[8902] = 8'hff ;
            rom[8903] = 8'he1 ;
            rom[8904] = 8'hf1 ;
            rom[8905] = 8'hf8 ;
            rom[8906] = 8'hfd ;
            rom[8907] = 8'h1e ;
            rom[8908] = 8'h04 ;
            rom[8909] = 8'hf9 ;
            rom[8910] = 8'h1c ;
            rom[8911] = 8'hf3 ;
            rom[8912] = 8'h18 ;
            rom[8913] = 8'hf9 ;
            rom[8914] = 8'h07 ;
            rom[8915] = 8'hca ;
            rom[8916] = 8'h10 ;
            rom[8917] = 8'h05 ;
            rom[8918] = 8'h03 ;
            rom[8919] = 8'h18 ;
            rom[8920] = 8'h09 ;
            rom[8921] = 8'he4 ;
            rom[8922] = 8'hfd ;
            rom[8923] = 8'he7 ;
            rom[8924] = 8'hf5 ;
            rom[8925] = 8'h03 ;
            rom[8926] = 8'h1c ;
            rom[8927] = 8'h0e ;
            rom[8928] = 8'h24 ;
            rom[8929] = 8'hf2 ;
            rom[8930] = 8'hfd ;
            rom[8931] = 8'hfe ;
            rom[8932] = 8'hd4 ;
            rom[8933] = 8'h1c ;
            rom[8934] = 8'he4 ;
            rom[8935] = 8'hf6 ;
            rom[8936] = 8'hdc ;
            rom[8937] = 8'hfe ;
            rom[8938] = 8'h0e ;
            rom[8939] = 8'hf2 ;
            rom[8940] = 8'h18 ;
            rom[8941] = 8'h05 ;
            rom[8942] = 8'hdc ;
            rom[8943] = 8'h2f ;
            rom[8944] = 8'h0a ;
            rom[8945] = 8'heb ;
            rom[8946] = 8'h00 ;
            rom[8947] = 8'h00 ;
            rom[8948] = 8'hf0 ;
            rom[8949] = 8'hf9 ;
            rom[8950] = 8'h1b ;
            rom[8951] = 8'h20 ;
            rom[8952] = 8'hf9 ;
            rom[8953] = 8'h0e ;
            rom[8954] = 8'hf8 ;
            rom[8955] = 8'h03 ;
            rom[8956] = 8'h00 ;
            rom[8957] = 8'h33 ;
            rom[8958] = 8'h06 ;
            rom[8959] = 8'h0b ;
            rom[8960] = 8'hf3 ;
            rom[8961] = 8'hfd ;
            rom[8962] = 8'h1e ;
            rom[8963] = 8'hde ;
            rom[8964] = 8'h05 ;
            rom[8965] = 8'h06 ;
            rom[8966] = 8'he2 ;
            rom[8967] = 8'h0a ;
            rom[8968] = 8'hfd ;
            rom[8969] = 8'h13 ;
            rom[8970] = 8'h03 ;
            rom[8971] = 8'hee ;
            rom[8972] = 8'h0c ;
            rom[8973] = 8'hee ;
            rom[8974] = 8'hfd ;
            rom[8975] = 8'h12 ;
            rom[8976] = 8'h0b ;
            rom[8977] = 8'hff ;
            rom[8978] = 8'he7 ;
            rom[8979] = 8'hfd ;
            rom[8980] = 8'hfb ;
            rom[8981] = 8'hef ;
            rom[8982] = 8'h11 ;
            rom[8983] = 8'hea ;
            rom[8984] = 8'ha2 ;
            rom[8985] = 8'hf7 ;
            rom[8986] = 8'hc1 ;
            rom[8987] = 8'h04 ;
            rom[8988] = 8'hc1 ;
            rom[8989] = 8'he3 ;
            rom[8990] = 8'h0a ;
            rom[8991] = 8'h04 ;
            rom[8992] = 8'h30 ;
            rom[8993] = 8'he6 ;
            rom[8994] = 8'h06 ;
            rom[8995] = 8'h18 ;
            rom[8996] = 8'he4 ;
            rom[8997] = 8'h03 ;
            rom[8998] = 8'he6 ;
            rom[8999] = 8'h12 ;
            rom[9000] = 8'h17 ;
            rom[9001] = 8'h01 ;
            rom[9002] = 8'hff ;
            rom[9003] = 8'h18 ;
            rom[9004] = 8'heb ;
            rom[9005] = 8'hd2 ;
            rom[9006] = 8'he6 ;
            rom[9007] = 8'h09 ;
            rom[9008] = 8'hf5 ;
            rom[9009] = 8'hed ;
            rom[9010] = 8'h02 ;
            rom[9011] = 8'he4 ;
            rom[9012] = 8'h10 ;
            rom[9013] = 8'he9 ;
            rom[9014] = 8'hff ;
            rom[9015] = 8'h0e ;
            rom[9016] = 8'h04 ;
            rom[9017] = 8'hd7 ;
            rom[9018] = 8'hd0 ;
            rom[9019] = 8'h06 ;
            rom[9020] = 8'hc3 ;
            rom[9021] = 8'hc0 ;
            rom[9022] = 8'h33 ;
            rom[9023] = 8'hf1 ;
            rom[9024] = 8'h0a ;
            rom[9025] = 8'h01 ;
            rom[9026] = 8'h1b ;
            rom[9027] = 8'hfc ;
            rom[9028] = 8'hda ;
            rom[9029] = 8'hf4 ;
            rom[9030] = 8'h1f ;
            rom[9031] = 8'hfc ;
            rom[9032] = 8'h00 ;
            rom[9033] = 8'hf1 ;
            rom[9034] = 8'hf1 ;
            rom[9035] = 8'hfb ;
            rom[9036] = 8'hae ;
            rom[9037] = 8'he2 ;
            rom[9038] = 8'h0a ;
            rom[9039] = 8'h10 ;
            rom[9040] = 8'hfe ;
            rom[9041] = 8'hf6 ;
            rom[9042] = 8'h0a ;
            rom[9043] = 8'hc7 ;
            rom[9044] = 8'hda ;
            rom[9045] = 8'h00 ;
            rom[9046] = 8'hfc ;
            rom[9047] = 8'h07 ;
            rom[9048] = 8'h11 ;
            rom[9049] = 8'h01 ;
            rom[9050] = 8'h13 ;
            rom[9051] = 8'he8 ;
            rom[9052] = 8'h18 ;
            rom[9053] = 8'heb ;
            rom[9054] = 8'h0b ;
            rom[9055] = 8'h09 ;
            rom[9056] = 8'h14 ;
            rom[9057] = 8'hf6 ;
            rom[9058] = 8'h05 ;
            rom[9059] = 8'h28 ;
            rom[9060] = 8'h00 ;
            rom[9061] = 8'h0b ;
            rom[9062] = 8'hdd ;
            rom[9063] = 8'h17 ;
            rom[9064] = 8'hea ;
            rom[9065] = 8'h0d ;
            rom[9066] = 8'h1c ;
            rom[9067] = 8'hee ;
            rom[9068] = 8'hc7 ;
            rom[9069] = 8'he6 ;
            rom[9070] = 8'hdb ;
            rom[9071] = 8'hcb ;
            rom[9072] = 8'hfa ;
            rom[9073] = 8'hfa ;
            rom[9074] = 8'h18 ;
            rom[9075] = 8'heb ;
            rom[9076] = 8'hd1 ;
            rom[9077] = 8'hf5 ;
            rom[9078] = 8'hd3 ;
            rom[9079] = 8'h16 ;
            rom[9080] = 8'h0a ;
            rom[9081] = 8'h0b ;
            rom[9082] = 8'h08 ;
            rom[9083] = 8'he5 ;
            rom[9084] = 8'h02 ;
            rom[9085] = 8'hff ;
            rom[9086] = 8'he2 ;
            rom[9087] = 8'h09 ;
            rom[9088] = 8'h29 ;
            rom[9089] = 8'h11 ;
            rom[9090] = 8'h07 ;
            rom[9091] = 8'hf6 ;
            rom[9092] = 8'he1 ;
            rom[9093] = 8'h0e ;
            rom[9094] = 8'hd9 ;
            rom[9095] = 8'hec ;
            rom[9096] = 8'h0f ;
            rom[9097] = 8'hf7 ;
            rom[9098] = 8'h05 ;
            rom[9099] = 8'h21 ;
            rom[9100] = 8'hdc ;
            rom[9101] = 8'hf3 ;
            rom[9102] = 8'h25 ;
            rom[9103] = 8'hf6 ;
            rom[9104] = 8'hf9 ;
            rom[9105] = 8'he2 ;
            rom[9106] = 8'h16 ;
            rom[9107] = 8'he6 ;
            rom[9108] = 8'hfe ;
            rom[9109] = 8'h05 ;
            rom[9110] = 8'he4 ;
            rom[9111] = 8'haa ;
            rom[9112] = 8'hf8 ;
            rom[9113] = 8'h15 ;
            rom[9114] = 8'hec ;
            rom[9115] = 8'h00 ;
            rom[9116] = 8'hfd ;
            rom[9117] = 8'h1c ;
            rom[9118] = 8'h04 ;
            rom[9119] = 8'hf0 ;
            rom[9120] = 8'h21 ;
            rom[9121] = 8'h17 ;
            rom[9122] = 8'h0e ;
            rom[9123] = 8'h1d ;
            rom[9124] = 8'he9 ;
            rom[9125] = 8'h11 ;
            rom[9126] = 8'hff ;
            rom[9127] = 8'h06 ;
            rom[9128] = 8'hf0 ;
            rom[9129] = 8'h19 ;
            rom[9130] = 8'hff ;
            rom[9131] = 8'h0c ;
            rom[9132] = 8'h08 ;
            rom[9133] = 8'hec ;
            rom[9134] = 8'h09 ;
            rom[9135] = 8'hee ;
            rom[9136] = 8'h1d ;
            rom[9137] = 8'h01 ;
            rom[9138] = 8'hf8 ;
            rom[9139] = 8'h18 ;
            rom[9140] = 8'h14 ;
            rom[9141] = 8'he4 ;
            rom[9142] = 8'hf7 ;
            rom[9143] = 8'he4 ;
            rom[9144] = 8'h13 ;
            rom[9145] = 8'hf7 ;
            rom[9146] = 8'hfb ;
            rom[9147] = 8'hed ;
            rom[9148] = 8'hf1 ;
            rom[9149] = 8'h02 ;
            rom[9150] = 8'h1a ;
            rom[9151] = 8'hf1 ;
            rom[9152] = 8'hf2 ;
            rom[9153] = 8'h01 ;
            rom[9154] = 8'h1d ;
            rom[9155] = 8'hfb ;
            rom[9156] = 8'hf8 ;
            rom[9157] = 8'h0c ;
            rom[9158] = 8'hf8 ;
            rom[9159] = 8'heb ;
            rom[9160] = 8'hfa ;
            rom[9161] = 8'h11 ;
            rom[9162] = 8'h05 ;
            rom[9163] = 8'h2c ;
            rom[9164] = 8'hf7 ;
            rom[9165] = 8'h01 ;
            rom[9166] = 8'h06 ;
            rom[9167] = 8'hf0 ;
            rom[9168] = 8'hfb ;
            rom[9169] = 8'ha8 ;
            rom[9170] = 8'hd8 ;
            rom[9171] = 8'hec ;
            rom[9172] = 8'hee ;
            rom[9173] = 8'hf1 ;
            rom[9174] = 8'he2 ;
            rom[9175] = 8'hfe ;
            rom[9176] = 8'hf6 ;
            rom[9177] = 8'hf9 ;
            rom[9178] = 8'hd4 ;
            rom[9179] = 8'h08 ;
            rom[9180] = 8'h12 ;
            rom[9181] = 8'hf1 ;
            rom[9182] = 8'h24 ;
            rom[9183] = 8'hea ;
            rom[9184] = 8'h17 ;
            rom[9185] = 8'h0c ;
            rom[9186] = 8'h09 ;
            rom[9187] = 8'hf8 ;
            rom[9188] = 8'hcf ;
            rom[9189] = 8'h1f ;
            rom[9190] = 8'he5 ;
            rom[9191] = 8'h12 ;
            rom[9192] = 8'h09 ;
            rom[9193] = 8'h06 ;
            rom[9194] = 8'hff ;
            rom[9195] = 8'h11 ;
            rom[9196] = 8'hed ;
            rom[9197] = 8'he4 ;
            rom[9198] = 8'he5 ;
            rom[9199] = 8'h1a ;
            rom[9200] = 8'he2 ;
            rom[9201] = 8'hfa ;
            rom[9202] = 8'h1e ;
            rom[9203] = 8'hfa ;
            rom[9204] = 8'hf0 ;
            rom[9205] = 8'hf2 ;
            rom[9206] = 8'h11 ;
            rom[9207] = 8'h12 ;
            rom[9208] = 8'hff ;
            rom[9209] = 8'hf0 ;
            rom[9210] = 8'hdd ;
            rom[9211] = 8'hd6 ;
            rom[9212] = 8'hc2 ;
            rom[9213] = 8'h10 ;
            rom[9214] = 8'h31 ;
            rom[9215] = 8'h08 ;
            rom[9216] = 8'h08 ;
            rom[9217] = 8'h11 ;
            rom[9218] = 8'hf6 ;
            rom[9219] = 8'h11 ;
            rom[9220] = 8'h03 ;
            rom[9221] = 8'he9 ;
            rom[9222] = 8'hf0 ;
            rom[9223] = 8'hef ;
            rom[9224] = 8'h09 ;
            rom[9225] = 8'hee ;
            rom[9226] = 8'hf9 ;
            rom[9227] = 8'hf1 ;
            rom[9228] = 8'h01 ;
            rom[9229] = 8'h09 ;
            rom[9230] = 8'he7 ;
            rom[9231] = 8'h18 ;
            rom[9232] = 8'h09 ;
            rom[9233] = 8'h0e ;
            rom[9234] = 8'hfa ;
            rom[9235] = 8'hed ;
            rom[9236] = 8'h03 ;
            rom[9237] = 8'h08 ;
            rom[9238] = 8'hf2 ;
            rom[9239] = 8'hdc ;
            rom[9240] = 8'hd8 ;
            rom[9241] = 8'hf1 ;
            rom[9242] = 8'hdd ;
            rom[9243] = 8'h08 ;
            rom[9244] = 8'hd2 ;
            rom[9245] = 8'h0b ;
            rom[9246] = 8'he5 ;
            rom[9247] = 8'h10 ;
            rom[9248] = 8'hf4 ;
            rom[9249] = 8'h10 ;
            rom[9250] = 8'h06 ;
            rom[9251] = 8'hc8 ;
            rom[9252] = 8'hec ;
            rom[9253] = 8'h18 ;
            rom[9254] = 8'h20 ;
            rom[9255] = 8'hed ;
            rom[9256] = 8'h12 ;
            rom[9257] = 8'h11 ;
            rom[9258] = 8'h12 ;
            rom[9259] = 8'hfc ;
            rom[9260] = 8'hf0 ;
            rom[9261] = 8'hc3 ;
            rom[9262] = 8'hf3 ;
            rom[9263] = 8'h0b ;
            rom[9264] = 8'hff ;
            rom[9265] = 8'hfe ;
            rom[9266] = 8'hec ;
            rom[9267] = 8'h05 ;
            rom[9268] = 8'hfd ;
            rom[9269] = 8'hb5 ;
            rom[9270] = 8'h0d ;
            rom[9271] = 8'h00 ;
            rom[9272] = 8'he2 ;
            rom[9273] = 8'hf7 ;
            rom[9274] = 8'hf2 ;
            rom[9275] = 8'h04 ;
            rom[9276] = 8'hd4 ;
            rom[9277] = 8'hde ;
            rom[9278] = 8'h17 ;
            rom[9279] = 8'hcf ;
            rom[9280] = 8'h0b ;
            rom[9281] = 8'hf9 ;
            rom[9282] = 8'h0a ;
            rom[9283] = 8'hd0 ;
            rom[9284] = 8'h19 ;
            rom[9285] = 8'h06 ;
            rom[9286] = 8'h0f ;
            rom[9287] = 8'h00 ;
            rom[9288] = 8'hfd ;
            rom[9289] = 8'h06 ;
            rom[9290] = 8'hde ;
            rom[9291] = 8'hb6 ;
            rom[9292] = 8'h01 ;
            rom[9293] = 8'hec ;
            rom[9294] = 8'he5 ;
            rom[9295] = 8'h02 ;
            rom[9296] = 8'h12 ;
            rom[9297] = 8'h0b ;
            rom[9298] = 8'h13 ;
            rom[9299] = 8'h02 ;
            rom[9300] = 8'h0a ;
            rom[9301] = 8'hfb ;
            rom[9302] = 8'h1c ;
            rom[9303] = 8'h14 ;
            rom[9304] = 8'hea ;
            rom[9305] = 8'h02 ;
            rom[9306] = 8'hf7 ;
            rom[9307] = 8'hd4 ;
            rom[9308] = 8'h0f ;
            rom[9309] = 8'h1e ;
            rom[9310] = 8'he2 ;
            rom[9311] = 8'hf5 ;
            rom[9312] = 8'h16 ;
            rom[9313] = 8'hf4 ;
            rom[9314] = 8'hf8 ;
            rom[9315] = 8'he6 ;
            rom[9316] = 8'h1e ;
            rom[9317] = 8'h18 ;
            rom[9318] = 8'h17 ;
            rom[9319] = 8'he8 ;
            rom[9320] = 8'h02 ;
            rom[9321] = 8'h01 ;
            rom[9322] = 8'hfe ;
            rom[9323] = 8'hd8 ;
            rom[9324] = 8'h02 ;
            rom[9325] = 8'h15 ;
            rom[9326] = 8'he7 ;
            rom[9327] = 8'h26 ;
            rom[9328] = 8'hf2 ;
            rom[9329] = 8'hf3 ;
            rom[9330] = 8'hff ;
            rom[9331] = 8'hd2 ;
            rom[9332] = 8'h09 ;
            rom[9333] = 8'h07 ;
            rom[9334] = 8'h07 ;
            rom[9335] = 8'h14 ;
            rom[9336] = 8'h01 ;
            rom[9337] = 8'h09 ;
            rom[9338] = 8'h0d ;
            rom[9339] = 8'h0b ;
            rom[9340] = 8'hf9 ;
            rom[9341] = 8'hec ;
            rom[9342] = 8'h1b ;
            rom[9343] = 8'he3 ;
            rom[9344] = 8'hf4 ;
            rom[9345] = 8'hfe ;
            rom[9346] = 8'h12 ;
            rom[9347] = 8'h05 ;
            rom[9348] = 8'h08 ;
            rom[9349] = 8'hff ;
            rom[9350] = 8'h1a ;
            rom[9351] = 8'h11 ;
            rom[9352] = 8'h1a ;
            rom[9353] = 8'hfb ;
            rom[9354] = 8'h0b ;
            rom[9355] = 8'hfd ;
            rom[9356] = 8'he0 ;
            rom[9357] = 8'hb3 ;
            rom[9358] = 8'hfc ;
            rom[9359] = 8'h07 ;
            rom[9360] = 8'hf9 ;
            rom[9361] = 8'h07 ;
            rom[9362] = 8'hf9 ;
            rom[9363] = 8'h14 ;
            rom[9364] = 8'hff ;
            rom[9365] = 8'hfd ;
            rom[9366] = 8'h19 ;
            rom[9367] = 8'h02 ;
            rom[9368] = 8'hbe ;
            rom[9369] = 8'hfd ;
            rom[9370] = 8'he0 ;
            rom[9371] = 8'h21 ;
            rom[9372] = 8'hc1 ;
            rom[9373] = 8'hf1 ;
            rom[9374] = 8'hf1 ;
            rom[9375] = 8'hf2 ;
            rom[9376] = 8'h06 ;
            rom[9377] = 8'hf5 ;
            rom[9378] = 8'hf5 ;
            rom[9379] = 8'hff ;
            rom[9380] = 8'h12 ;
            rom[9381] = 8'h12 ;
            rom[9382] = 8'hfa ;
            rom[9383] = 8'h0c ;
            rom[9384] = 8'h17 ;
            rom[9385] = 8'h06 ;
            rom[9386] = 8'h0b ;
            rom[9387] = 8'h26 ;
            rom[9388] = 8'hf0 ;
            rom[9389] = 8'hb5 ;
            rom[9390] = 8'h05 ;
            rom[9391] = 8'h02 ;
            rom[9392] = 8'hdf ;
            rom[9393] = 8'h0b ;
            rom[9394] = 8'hee ;
            rom[9395] = 8'hfa ;
            rom[9396] = 8'h01 ;
            rom[9397] = 8'hd3 ;
            rom[9398] = 8'hf4 ;
            rom[9399] = 8'hfd ;
            rom[9400] = 8'h08 ;
            rom[9401] = 8'hd9 ;
            rom[9402] = 8'h14 ;
            rom[9403] = 8'h0e ;
            rom[9404] = 8'hd9 ;
            rom[9405] = 8'heb ;
            rom[9406] = 8'hf8 ;
            rom[9407] = 8'hc8 ;
            rom[9408] = 8'hea ;
            rom[9409] = 8'h00 ;
            rom[9410] = 8'hef ;
            rom[9411] = 8'h0c ;
            rom[9412] = 8'hf4 ;
            rom[9413] = 8'hb9 ;
            rom[9414] = 8'h00 ;
            rom[9415] = 8'hf1 ;
            rom[9416] = 8'h03 ;
            rom[9417] = 8'hcc ;
            rom[9418] = 8'hba ;
            rom[9419] = 8'h03 ;
            rom[9420] = 8'hda ;
            rom[9421] = 8'hdf ;
            rom[9422] = 8'h01 ;
            rom[9423] = 8'h06 ;
            rom[9424] = 8'h10 ;
            rom[9425] = 8'h08 ;
            rom[9426] = 8'h0d ;
            rom[9427] = 8'hfc ;
            rom[9428] = 8'hfd ;
            rom[9429] = 8'h15 ;
            rom[9430] = 8'hea ;
            rom[9431] = 8'hff ;
            rom[9432] = 8'h03 ;
            rom[9433] = 8'h02 ;
            rom[9434] = 8'h2c ;
            rom[9435] = 8'he1 ;
            rom[9436] = 8'h16 ;
            rom[9437] = 8'h0e ;
            rom[9438] = 8'h07 ;
            rom[9439] = 8'hd8 ;
            rom[9440] = 8'h06 ;
            rom[9441] = 8'he6 ;
            rom[9442] = 8'hf8 ;
            rom[9443] = 8'he3 ;
            rom[9444] = 8'hf5 ;
            rom[9445] = 8'h10 ;
            rom[9446] = 8'hf0 ;
            rom[9447] = 8'h06 ;
            rom[9448] = 8'h0d ;
            rom[9449] = 8'hb6 ;
            rom[9450] = 8'he3 ;
            rom[9451] = 8'hf8 ;
            rom[9452] = 8'hfd ;
            rom[9453] = 8'h0c ;
            rom[9454] = 8'hdb ;
            rom[9455] = 8'h15 ;
            rom[9456] = 8'h01 ;
            rom[9457] = 8'hcf ;
            rom[9458] = 8'h0c ;
            rom[9459] = 8'h0b ;
            rom[9460] = 8'hfc ;
            rom[9461] = 8'h09 ;
            rom[9462] = 8'had ;
            rom[9463] = 8'hfd ;
            rom[9464] = 8'hea ;
            rom[9465] = 8'h14 ;
            rom[9466] = 8'h03 ;
            rom[9467] = 8'h03 ;
            rom[9468] = 8'hfa ;
            rom[9469] = 8'h0c ;
            rom[9470] = 8'h10 ;
            rom[9471] = 8'h0b ;
            rom[9472] = 8'h1f ;
            rom[9473] = 8'h06 ;
            rom[9474] = 8'hdb ;
            rom[9475] = 8'hea ;
            rom[9476] = 8'h03 ;
            rom[9477] = 8'h1b ;
            rom[9478] = 8'h13 ;
            rom[9479] = 8'h04 ;
            rom[9480] = 8'h03 ;
            rom[9481] = 8'hfd ;
            rom[9482] = 8'h09 ;
            rom[9483] = 8'hea ;
            rom[9484] = 8'h13 ;
            rom[9485] = 8'hee ;
            rom[9486] = 8'hce ;
            rom[9487] = 8'h02 ;
            rom[9488] = 8'h13 ;
            rom[9489] = 8'h0f ;
            rom[9490] = 8'h1d ;
            rom[9491] = 8'h0c ;
            rom[9492] = 8'he0 ;
            rom[9493] = 8'hf8 ;
            rom[9494] = 8'h08 ;
            rom[9495] = 8'h08 ;
            rom[9496] = 8'hcd ;
            rom[9497] = 8'hed ;
            rom[9498] = 8'hdf ;
            rom[9499] = 8'hd9 ;
            rom[9500] = 8'hf2 ;
            rom[9501] = 8'h07 ;
            rom[9502] = 8'hd6 ;
            rom[9503] = 8'hfc ;
            rom[9504] = 8'hfa ;
            rom[9505] = 8'h05 ;
            rom[9506] = 8'h14 ;
            rom[9507] = 8'hd2 ;
            rom[9508] = 8'h12 ;
            rom[9509] = 8'h0f ;
            rom[9510] = 8'hf7 ;
            rom[9511] = 8'hf3 ;
            rom[9512] = 8'h09 ;
            rom[9513] = 8'hef ;
            rom[9514] = 8'h09 ;
            rom[9515] = 8'hee ;
            rom[9516] = 8'hda ;
            rom[9517] = 8'hf7 ;
            rom[9518] = 8'h07 ;
            rom[9519] = 8'hf4 ;
            rom[9520] = 8'hfd ;
            rom[9521] = 8'hf3 ;
            rom[9522] = 8'hd9 ;
            rom[9523] = 8'h1d ;
            rom[9524] = 8'h00 ;
            rom[9525] = 8'hda ;
            rom[9526] = 8'h07 ;
            rom[9527] = 8'hf5 ;
            rom[9528] = 8'h01 ;
            rom[9529] = 8'haf ;
            rom[9530] = 8'h03 ;
            rom[9531] = 8'h15 ;
            rom[9532] = 8'hf3 ;
            rom[9533] = 8'he3 ;
            rom[9534] = 8'heb ;
            rom[9535] = 8'hdb ;
            rom[9536] = 8'h16 ;
            rom[9537] = 8'h06 ;
            rom[9538] = 8'h04 ;
            rom[9539] = 8'h0a ;
            rom[9540] = 8'h04 ;
            rom[9541] = 8'hb6 ;
            rom[9542] = 8'hde ;
            rom[9543] = 8'hfc ;
            rom[9544] = 8'h16 ;
            rom[9545] = 8'hc9 ;
            rom[9546] = 8'h08 ;
            rom[9547] = 8'h25 ;
            rom[9548] = 8'h10 ;
            rom[9549] = 8'hf9 ;
            rom[9550] = 8'hf8 ;
            rom[9551] = 8'h14 ;
            rom[9552] = 8'h15 ;
            rom[9553] = 8'h10 ;
            rom[9554] = 8'h18 ;
            rom[9555] = 8'h11 ;
            rom[9556] = 8'hfd ;
            rom[9557] = 8'h02 ;
            rom[9558] = 8'hff ;
            rom[9559] = 8'hf2 ;
            rom[9560] = 8'h14 ;
            rom[9561] = 8'hf8 ;
            rom[9562] = 8'he1 ;
            rom[9563] = 8'hf0 ;
            rom[9564] = 8'hfd ;
            rom[9565] = 8'h05 ;
            rom[9566] = 8'hf0 ;
            rom[9567] = 8'h10 ;
            rom[9568] = 8'h16 ;
            rom[9569] = 8'hfe ;
            rom[9570] = 8'hde ;
            rom[9571] = 8'heb ;
            rom[9572] = 8'he0 ;
            rom[9573] = 8'heb ;
            rom[9574] = 8'hed ;
            rom[9575] = 8'hf7 ;
            rom[9576] = 8'hd6 ;
            rom[9577] = 8'h08 ;
            rom[9578] = 8'h0a ;
            rom[9579] = 8'hf8 ;
            rom[9580] = 8'h01 ;
            rom[9581] = 8'he2 ;
            rom[9582] = 8'hfe ;
            rom[9583] = 8'h0b ;
            rom[9584] = 8'h14 ;
            rom[9585] = 8'h02 ;
            rom[9586] = 8'hea ;
            rom[9587] = 8'h02 ;
            rom[9588] = 8'hd2 ;
            rom[9589] = 8'hec ;
            rom[9590] = 8'h13 ;
            rom[9591] = 8'hf7 ;
            rom[9592] = 8'hde ;
            rom[9593] = 8'hd0 ;
            rom[9594] = 8'h0b ;
            rom[9595] = 8'h19 ;
            rom[9596] = 8'hff ;
            rom[9597] = 8'hf5 ;
            rom[9598] = 8'h19 ;
            rom[9599] = 8'hf0 ;
            rom[9600] = 8'h12 ;
            rom[9601] = 8'hdc ;
            rom[9602] = 8'hfc ;
            rom[9603] = 8'he2 ;
            rom[9604] = 8'hd5 ;
            rom[9605] = 8'h07 ;
            rom[9606] = 8'hff ;
            rom[9607] = 8'he6 ;
            rom[9608] = 8'hf8 ;
            rom[9609] = 8'hf4 ;
            rom[9610] = 8'h09 ;
            rom[9611] = 8'h12 ;
            rom[9612] = 8'h0f ;
            rom[9613] = 8'hd3 ;
            rom[9614] = 8'hcd ;
            rom[9615] = 8'heb ;
            rom[9616] = 8'hf9 ;
            rom[9617] = 8'h12 ;
            rom[9618] = 8'hfa ;
            rom[9619] = 8'hd6 ;
            rom[9620] = 8'h00 ;
            rom[9621] = 8'he8 ;
            rom[9622] = 8'h14 ;
            rom[9623] = 8'h02 ;
            rom[9624] = 8'h10 ;
            rom[9625] = 8'hf2 ;
            rom[9626] = 8'hf5 ;
            rom[9627] = 8'hfe ;
            rom[9628] = 8'hf8 ;
            rom[9629] = 8'h21 ;
            rom[9630] = 8'he6 ;
            rom[9631] = 8'h0a ;
            rom[9632] = 8'h29 ;
            rom[9633] = 8'h0f ;
            rom[9634] = 8'hcd ;
            rom[9635] = 8'h09 ;
            rom[9636] = 8'h04 ;
            rom[9637] = 8'h13 ;
            rom[9638] = 8'hfb ;
            rom[9639] = 8'h1c ;
            rom[9640] = 8'heb ;
            rom[9641] = 8'hf6 ;
            rom[9642] = 8'h07 ;
            rom[9643] = 8'hea ;
            rom[9644] = 8'he8 ;
            rom[9645] = 8'hfb ;
            rom[9646] = 8'h13 ;
            rom[9647] = 8'hc6 ;
            rom[9648] = 8'hf1 ;
            rom[9649] = 8'hc5 ;
            rom[9650] = 8'hcf ;
            rom[9651] = 8'h0f ;
            rom[9652] = 8'hb7 ;
            rom[9653] = 8'hfd ;
            rom[9654] = 8'hf0 ;
            rom[9655] = 8'h0b ;
            rom[9656] = 8'h14 ;
            rom[9657] = 8'h0d ;
            rom[9658] = 8'hf4 ;
            rom[9659] = 8'h0e ;
            rom[9660] = 8'h10 ;
            rom[9661] = 8'hf9 ;
            rom[9662] = 8'h06 ;
            rom[9663] = 8'h07 ;
            rom[9664] = 8'h13 ;
            rom[9665] = 8'hfc ;
            rom[9666] = 8'h06 ;
            rom[9667] = 8'h07 ;
            rom[9668] = 8'he9 ;
            rom[9669] = 8'hf2 ;
            rom[9670] = 8'hef ;
            rom[9671] = 8'h0f ;
            rom[9672] = 8'h08 ;
            rom[9673] = 8'heb ;
            rom[9674] = 8'h00 ;
            rom[9675] = 8'h2e ;
            rom[9676] = 8'hf6 ;
            rom[9677] = 8'hf4 ;
            rom[9678] = 8'h0b ;
            rom[9679] = 8'hf4 ;
            rom[9680] = 8'hfe ;
            rom[9681] = 8'h00 ;
            rom[9682] = 8'h07 ;
            rom[9683] = 8'h20 ;
            rom[9684] = 8'hd2 ;
            rom[9685] = 8'h03 ;
            rom[9686] = 8'h08 ;
            rom[9687] = 8'hf4 ;
            rom[9688] = 8'h07 ;
            rom[9689] = 8'hfc ;
            rom[9690] = 8'hdd ;
            rom[9691] = 8'h0f ;
            rom[9692] = 8'hb9 ;
            rom[9693] = 8'he7 ;
            rom[9694] = 8'hec ;
            rom[9695] = 8'h06 ;
            rom[9696] = 8'hf1 ;
            rom[9697] = 8'he9 ;
            rom[9698] = 8'he2 ;
            rom[9699] = 8'hfc ;
            rom[9700] = 8'hed ;
            rom[9701] = 8'hf2 ;
            rom[9702] = 8'hfc ;
            rom[9703] = 8'he5 ;
            rom[9704] = 8'hf0 ;
            rom[9705] = 8'h13 ;
            rom[9706] = 8'h12 ;
            rom[9707] = 8'h10 ;
            rom[9708] = 8'h05 ;
            rom[9709] = 8'he2 ;
            rom[9710] = 8'h14 ;
            rom[9711] = 8'h19 ;
            rom[9712] = 8'hf4 ;
            rom[9713] = 8'h07 ;
            rom[9714] = 8'h11 ;
            rom[9715] = 8'h0f ;
            rom[9716] = 8'hd7 ;
            rom[9717] = 8'hf5 ;
            rom[9718] = 8'hf2 ;
            rom[9719] = 8'hf5 ;
            rom[9720] = 8'hdb ;
            rom[9721] = 8'hdb ;
            rom[9722] = 8'hfb ;
            rom[9723] = 8'h25 ;
            rom[9724] = 8'h17 ;
            rom[9725] = 8'h03 ;
            rom[9726] = 8'h0e ;
            rom[9727] = 8'hef ;
            rom[9728] = 8'h01 ;
            rom[9729] = 8'he1 ;
            rom[9730] = 8'h1b ;
            rom[9731] = 8'hc9 ;
            rom[9732] = 8'hff ;
            rom[9733] = 8'h05 ;
            rom[9734] = 8'h1a ;
            rom[9735] = 8'he9 ;
            rom[9736] = 8'hf8 ;
            rom[9737] = 8'he9 ;
            rom[9738] = 8'hfd ;
            rom[9739] = 8'hd4 ;
            rom[9740] = 8'h02 ;
            rom[9741] = 8'he6 ;
            rom[9742] = 8'hd0 ;
            rom[9743] = 8'hfd ;
            rom[9744] = 8'hf7 ;
            rom[9745] = 8'h06 ;
            rom[9746] = 8'hf4 ;
            rom[9747] = 8'h11 ;
            rom[9748] = 8'hd8 ;
            rom[9749] = 8'h09 ;
            rom[9750] = 8'hfb ;
            rom[9751] = 8'hea ;
            rom[9752] = 8'hda ;
            rom[9753] = 8'hee ;
            rom[9754] = 8'hd0 ;
            rom[9755] = 8'hfb ;
            rom[9756] = 8'hf7 ;
            rom[9757] = 8'hff ;
            rom[9758] = 8'hf6 ;
            rom[9759] = 8'he5 ;
            rom[9760] = 8'h20 ;
            rom[9761] = 8'hd3 ;
            rom[9762] = 8'hd8 ;
            rom[9763] = 8'h0e ;
            rom[9764] = 8'h21 ;
            rom[9765] = 8'h1f ;
            rom[9766] = 8'h00 ;
            rom[9767] = 8'h18 ;
            rom[9768] = 8'hf2 ;
            rom[9769] = 8'hee ;
            rom[9770] = 8'h1c ;
            rom[9771] = 8'hf5 ;
            rom[9772] = 8'hf6 ;
            rom[9773] = 8'hef ;
            rom[9774] = 8'he2 ;
            rom[9775] = 8'h0b ;
            rom[9776] = 8'hfd ;
            rom[9777] = 8'hd6 ;
            rom[9778] = 8'h09 ;
            rom[9779] = 8'hd3 ;
            rom[9780] = 8'he5 ;
            rom[9781] = 8'hfd ;
            rom[9782] = 8'hed ;
            rom[9783] = 8'h05 ;
            rom[9784] = 8'h1b ;
            rom[9785] = 8'hdd ;
            rom[9786] = 8'h00 ;
            rom[9787] = 8'hff ;
            rom[9788] = 8'h0c ;
            rom[9789] = 8'he8 ;
            rom[9790] = 8'h04 ;
            rom[9791] = 8'hff ;
            rom[9792] = 8'hf8 ;
            rom[9793] = 8'h26 ;
            rom[9794] = 8'hf8 ;
            rom[9795] = 8'hef ;
            rom[9796] = 8'he8 ;
            rom[9797] = 8'he1 ;
            rom[9798] = 8'h00 ;
            rom[9799] = 8'hf8 ;
            rom[9800] = 8'hf7 ;
            rom[9801] = 8'hed ;
            rom[9802] = 8'ha2 ;
            rom[9803] = 8'h0f ;
            rom[9804] = 8'he7 ;
            rom[9805] = 8'he1 ;
            rom[9806] = 8'hec ;
            rom[9807] = 8'h03 ;
            rom[9808] = 8'h0f ;
            rom[9809] = 8'h0c ;
            rom[9810] = 8'h0c ;
            rom[9811] = 8'hfe ;
            rom[9812] = 8'hd5 ;
            rom[9813] = 8'h0a ;
            rom[9814] = 8'hd3 ;
            rom[9815] = 8'h0b ;
            rom[9816] = 8'h0a ;
            rom[9817] = 8'hed ;
            rom[9818] = 8'h1f ;
            rom[9819] = 8'hdc ;
            rom[9820] = 8'hf1 ;
            rom[9821] = 8'h0d ;
            rom[9822] = 8'h16 ;
            rom[9823] = 8'he1 ;
            rom[9824] = 8'h18 ;
            rom[9825] = 8'he7 ;
            rom[9826] = 8'hf2 ;
            rom[9827] = 8'hd3 ;
            rom[9828] = 8'he4 ;
            rom[9829] = 8'h04 ;
            rom[9830] = 8'hfc ;
            rom[9831] = 8'h01 ;
            rom[9832] = 8'hfe ;
            rom[9833] = 8'hcc ;
            rom[9834] = 8'hf3 ;
            rom[9835] = 8'hf1 ;
            rom[9836] = 8'h0c ;
            rom[9837] = 8'h07 ;
            rom[9838] = 8'he1 ;
            rom[9839] = 8'h13 ;
            rom[9840] = 8'h14 ;
            rom[9841] = 8'hce ;
            rom[9842] = 8'hf4 ;
            rom[9843] = 8'h07 ;
            rom[9844] = 8'he2 ;
            rom[9845] = 8'h04 ;
            rom[9846] = 8'hc5 ;
            rom[9847] = 8'hfa ;
            rom[9848] = 8'hf1 ;
            rom[9849] = 8'h0f ;
            rom[9850] = 8'h02 ;
            rom[9851] = 8'h00 ;
            rom[9852] = 8'hfb ;
            rom[9853] = 8'h16 ;
            rom[9854] = 8'h09 ;
            rom[9855] = 8'hec ;
            rom[9856] = 8'hef ;
            rom[9857] = 8'h0f ;
            rom[9858] = 8'h07 ;
            rom[9859] = 8'hd3 ;
            rom[9860] = 8'heb ;
            rom[9861] = 8'he5 ;
            rom[9862] = 8'hf4 ;
            rom[9863] = 8'h0b ;
            rom[9864] = 8'hf2 ;
            rom[9865] = 8'hd0 ;
            rom[9866] = 8'he7 ;
            rom[9867] = 8'h06 ;
            rom[9868] = 8'h04 ;
            rom[9869] = 8'hf6 ;
            rom[9870] = 8'h09 ;
            rom[9871] = 8'h11 ;
            rom[9872] = 8'hfc ;
            rom[9873] = 8'h07 ;
            rom[9874] = 8'h19 ;
            rom[9875] = 8'hc7 ;
            rom[9876] = 8'hb3 ;
            rom[9877] = 8'hf1 ;
            rom[9878] = 8'h08 ;
            rom[9879] = 8'h20 ;
            rom[9880] = 8'h0f ;
            rom[9881] = 8'hdc ;
            rom[9882] = 8'h13 ;
            rom[9883] = 8'hbc ;
            rom[9884] = 8'hff ;
            rom[9885] = 8'h06 ;
            rom[9886] = 8'h02 ;
            rom[9887] = 8'h03 ;
            rom[9888] = 8'h1d ;
            rom[9889] = 8'hdc ;
            rom[9890] = 8'hd8 ;
            rom[9891] = 8'hcd ;
            rom[9892] = 8'hec ;
            rom[9893] = 8'h13 ;
            rom[9894] = 8'hff ;
            rom[9895] = 8'h19 ;
            rom[9896] = 8'hed ;
            rom[9897] = 8'hcf ;
            rom[9898] = 8'hf3 ;
            rom[9899] = 8'he2 ;
            rom[9900] = 8'h03 ;
            rom[9901] = 8'hf7 ;
            rom[9902] = 8'hfa ;
            rom[9903] = 8'hee ;
            rom[9904] = 8'h13 ;
            rom[9905] = 8'hc9 ;
            rom[9906] = 8'hf6 ;
            rom[9907] = 8'hf1 ;
            rom[9908] = 8'hb6 ;
            rom[9909] = 8'h02 ;
            rom[9910] = 8'hfa ;
            rom[9911] = 8'h0e ;
            rom[9912] = 8'h0d ;
            rom[9913] = 8'h08 ;
            rom[9914] = 8'h10 ;
            rom[9915] = 8'h01 ;
            rom[9916] = 8'h0d ;
            rom[9917] = 8'hfc ;
            rom[9918] = 8'hff ;
            rom[9919] = 8'h13 ;
            rom[9920] = 8'h01 ;
            rom[9921] = 8'h05 ;
            rom[9922] = 8'h06 ;
            rom[9923] = 8'hf6 ;
            rom[9924] = 8'hee ;
            rom[9925] = 8'hb2 ;
            rom[9926] = 8'hf0 ;
            rom[9927] = 8'h0d ;
            rom[9928] = 8'h12 ;
            rom[9929] = 8'hb9 ;
            rom[9930] = 8'he7 ;
            rom[9931] = 8'h16 ;
            rom[9932] = 8'he9 ;
            rom[9933] = 8'hd1 ;
            rom[9934] = 8'h07 ;
            rom[9935] = 8'h0e ;
            rom[9936] = 8'h0e ;
            rom[9937] = 8'h00 ;
            rom[9938] = 8'h1f ;
            rom[9939] = 8'h0e ;
            rom[9940] = 8'hd6 ;
            rom[9941] = 8'hfb ;
            rom[9942] = 8'h1f ;
            rom[9943] = 8'hfa ;
            rom[9944] = 8'h1d ;
            rom[9945] = 8'h12 ;
            rom[9946] = 8'h21 ;
            rom[9947] = 8'hef ;
            rom[9948] = 8'hf8 ;
            rom[9949] = 8'hd9 ;
            rom[9950] = 8'hf5 ;
            rom[9951] = 8'h03 ;
            rom[9952] = 8'h10 ;
            rom[9953] = 8'h00 ;
            rom[9954] = 8'hb0 ;
            rom[9955] = 8'hdc ;
            rom[9956] = 8'he9 ;
            rom[9957] = 8'h10 ;
            rom[9958] = 8'hfa ;
            rom[9959] = 8'hfb ;
            rom[9960] = 8'heb ;
            rom[9961] = 8'hfe ;
            rom[9962] = 8'h03 ;
            rom[9963] = 8'he2 ;
            rom[9964] = 8'hf1 ;
            rom[9965] = 8'h01 ;
            rom[9966] = 8'h04 ;
            rom[9967] = 8'h0b ;
            rom[9968] = 8'h08 ;
            rom[9969] = 8'h03 ;
            rom[9970] = 8'hf8 ;
            rom[9971] = 8'heb ;
            rom[9972] = 8'hdf ;
            rom[9973] = 8'hf2 ;
            rom[9974] = 8'hdc ;
            rom[9975] = 8'hf6 ;
            rom[9976] = 8'he5 ;
            rom[9977] = 8'h17 ;
            rom[9978] = 8'h07 ;
            rom[9979] = 8'hfb ;
            rom[9980] = 8'h03 ;
            rom[9981] = 8'h01 ;
            rom[9982] = 8'hfe ;
            rom[9983] = 8'h06 ;
            rom[9984] = 8'h1b ;
            rom[9985] = 8'h05 ;
            rom[9986] = 8'hee ;
            rom[9987] = 8'h0c ;
            rom[9988] = 8'hec ;
            rom[9989] = 8'hdf ;
            rom[9990] = 8'hed ;
            rom[9991] = 8'h14 ;
            rom[9992] = 8'h19 ;
            rom[9993] = 8'hcb ;
            rom[9994] = 8'h14 ;
            rom[9995] = 8'h12 ;
            rom[9996] = 8'hf7 ;
            rom[9997] = 8'hfd ;
            rom[9998] = 8'he8 ;
            rom[9999] = 8'hfa ;
            rom[10000] = 8'h19 ;
            rom[10001] = 8'h2d ;
            rom[10002] = 8'h1c ;
            rom[10003] = 8'h01 ;
            rom[10004] = 8'he6 ;
            rom[10005] = 8'h0d ;
            rom[10006] = 8'hfe ;
            rom[10007] = 8'hf0 ;
            rom[10008] = 8'hf0 ;
            rom[10009] = 8'hf8 ;
            rom[10010] = 8'he2 ;
            rom[10011] = 8'hf3 ;
            rom[10012] = 8'he6 ;
            rom[10013] = 8'hea ;
            rom[10014] = 8'he6 ;
            rom[10015] = 8'h11 ;
            rom[10016] = 8'he4 ;
            rom[10017] = 8'h03 ;
            rom[10018] = 8'heb ;
            rom[10019] = 8'h03 ;
            rom[10020] = 8'he4 ;
            rom[10021] = 8'heb ;
            rom[10022] = 8'h0e ;
            rom[10023] = 8'hf8 ;
            rom[10024] = 8'hec ;
            rom[10025] = 8'h06 ;
            rom[10026] = 8'h09 ;
            rom[10027] = 8'hf8 ;
            rom[10028] = 8'hfe ;
            rom[10029] = 8'hfb ;
            rom[10030] = 8'h12 ;
            rom[10031] = 8'h04 ;
            rom[10032] = 8'h02 ;
            rom[10033] = 8'hf8 ;
            rom[10034] = 8'hde ;
            rom[10035] = 8'hed ;
            rom[10036] = 8'h03 ;
            rom[10037] = 8'he1 ;
            rom[10038] = 8'hfe ;
            rom[10039] = 8'h0f ;
            rom[10040] = 8'hbe ;
            rom[10041] = 8'hd2 ;
            rom[10042] = 8'h25 ;
            rom[10043] = 8'h10 ;
            rom[10044] = 8'he3 ;
            rom[10045] = 8'hf7 ;
            rom[10046] = 8'h11 ;
            rom[10047] = 8'h07 ;
            rom[10048] = 8'h0f ;
            rom[10049] = 8'h0b ;
            rom[10050] = 8'he2 ;
            rom[10051] = 8'hd8 ;
            rom[10052] = 8'h1d ;
            rom[10053] = 8'h19 ;
            rom[10054] = 8'h12 ;
            rom[10055] = 8'hc7 ;
            rom[10056] = 8'hfd ;
            rom[10057] = 8'hff ;
            rom[10058] = 8'h06 ;
            rom[10059] = 8'hfc ;
            rom[10060] = 8'h02 ;
            rom[10061] = 8'hee ;
            rom[10062] = 8'h09 ;
            rom[10063] = 8'hdc ;
            rom[10064] = 8'h0b ;
            rom[10065] = 8'h0e ;
            rom[10066] = 8'h02 ;
            rom[10067] = 8'he2 ;
            rom[10068] = 8'hcb ;
            rom[10069] = 8'hc4 ;
            rom[10070] = 8'hf5 ;
            rom[10071] = 8'h00 ;
            rom[10072] = 8'h07 ;
            rom[10073] = 8'hf9 ;
            rom[10074] = 8'h0f ;
            rom[10075] = 8'he0 ;
            rom[10076] = 8'hfb ;
            rom[10077] = 8'hf8 ;
            rom[10078] = 8'hf5 ;
            rom[10079] = 8'h0b ;
            rom[10080] = 8'h04 ;
            rom[10081] = 8'hed ;
            rom[10082] = 8'h01 ;
            rom[10083] = 8'hfa ;
            rom[10084] = 8'h13 ;
            rom[10085] = 8'h0a ;
            rom[10086] = 8'h09 ;
            rom[10087] = 8'hfd ;
            rom[10088] = 8'hf3 ;
            rom[10089] = 8'hd7 ;
            rom[10090] = 8'h03 ;
            rom[10091] = 8'hf1 ;
            rom[10092] = 8'hfb ;
            rom[10093] = 8'hf9 ;
            rom[10094] = 8'hd9 ;
            rom[10095] = 8'hf1 ;
            rom[10096] = 8'h00 ;
            rom[10097] = 8'hd9 ;
            rom[10098] = 8'h0a ;
            rom[10099] = 8'h03 ;
            rom[10100] = 8'hbf ;
            rom[10101] = 8'h09 ;
            rom[10102] = 8'h19 ;
            rom[10103] = 8'hfc ;
            rom[10104] = 8'hfd ;
            rom[10105] = 8'h2b ;
            rom[10106] = 8'he4 ;
            rom[10107] = 8'h0f ;
            rom[10108] = 8'h04 ;
            rom[10109] = 8'hfb ;
            rom[10110] = 8'hfb ;
            rom[10111] = 8'h03 ;
            rom[10112] = 8'h0a ;
            rom[10113] = 8'h08 ;
            rom[10114] = 8'h0a ;
            rom[10115] = 8'hcc ;
            rom[10116] = 8'hec ;
            rom[10117] = 8'hfc ;
            rom[10118] = 8'hf0 ;
            rom[10119] = 8'hbe ;
            rom[10120] = 8'hf6 ;
            rom[10121] = 8'h21 ;
            rom[10122] = 8'h0d ;
            rom[10123] = 8'h02 ;
            rom[10124] = 8'hfc ;
            rom[10125] = 8'h03 ;
            rom[10126] = 8'hf6 ;
            rom[10127] = 8'hfc ;
            rom[10128] = 8'h00 ;
            rom[10129] = 8'h19 ;
            rom[10130] = 8'hdc ;
            rom[10131] = 8'h14 ;
            rom[10132] = 8'hf9 ;
            rom[10133] = 8'hf3 ;
            rom[10134] = 8'he5 ;
            rom[10135] = 8'hdd ;
            rom[10136] = 8'hbf ;
            rom[10137] = 8'he5 ;
            rom[10138] = 8'he3 ;
            rom[10139] = 8'h1e ;
            rom[10140] = 8'hfb ;
            rom[10141] = 8'h08 ;
            rom[10142] = 8'h09 ;
            rom[10143] = 8'hfe ;
            rom[10144] = 8'heb ;
            rom[10145] = 8'h07 ;
            rom[10146] = 8'hee ;
            rom[10147] = 8'h16 ;
            rom[10148] = 8'hf8 ;
            rom[10149] = 8'h1a ;
            rom[10150] = 8'hf5 ;
            rom[10151] = 8'h03 ;
            rom[10152] = 8'hf7 ;
            rom[10153] = 8'hfb ;
            rom[10154] = 8'hde ;
            rom[10155] = 8'h07 ;
            rom[10156] = 8'h13 ;
            rom[10157] = 8'hf1 ;
            rom[10158] = 8'hfa ;
            rom[10159] = 8'hd6 ;
            rom[10160] = 8'h1f ;
            rom[10161] = 8'hdb ;
            rom[10162] = 8'hf8 ;
            rom[10163] = 8'hc7 ;
            rom[10164] = 8'h14 ;
            rom[10165] = 8'hf5 ;
            rom[10166] = 8'hf0 ;
            rom[10167] = 8'h20 ;
            rom[10168] = 8'h03 ;
            rom[10169] = 8'h0f ;
            rom[10170] = 8'he1 ;
            rom[10171] = 8'he3 ;
            rom[10172] = 8'hf7 ;
            rom[10173] = 8'he1 ;
            rom[10174] = 8'h12 ;
            rom[10175] = 8'h14 ;
            rom[10176] = 8'h07 ;
            rom[10177] = 8'hf8 ;
            rom[10178] = 8'hea ;
            rom[10179] = 8'h1f ;
            rom[10180] = 8'h1b ;
            rom[10181] = 8'h11 ;
            rom[10182] = 8'h00 ;
            rom[10183] = 8'h03 ;
            rom[10184] = 8'h15 ;
            rom[10185] = 8'hf6 ;
            rom[10186] = 8'h1b ;
            rom[10187] = 8'h02 ;
            rom[10188] = 8'h13 ;
            rom[10189] = 8'hfe ;
            rom[10190] = 8'h08 ;
            rom[10191] = 8'hf0 ;
            rom[10192] = 8'h0a ;
            rom[10193] = 8'h09 ;
            rom[10194] = 8'hfa ;
            rom[10195] = 8'hd4 ;
            rom[10196] = 8'hf9 ;
            rom[10197] = 8'hf1 ;
            rom[10198] = 8'h0b ;
            rom[10199] = 8'h0a ;
            rom[10200] = 8'h03 ;
            rom[10201] = 8'h0d ;
            rom[10202] = 8'h05 ;
            rom[10203] = 8'h0b ;
            rom[10204] = 8'hf5 ;
            rom[10205] = 8'hfa ;
            rom[10206] = 8'h05 ;
            rom[10207] = 8'hfc ;
            rom[10208] = 8'h0c ;
            rom[10209] = 8'he3 ;
            rom[10210] = 8'hf9 ;
            rom[10211] = 8'h08 ;
            rom[10212] = 8'h23 ;
            rom[10213] = 8'h13 ;
            rom[10214] = 8'h07 ;
            rom[10215] = 8'he0 ;
            rom[10216] = 8'hd2 ;
            rom[10217] = 8'hdc ;
            rom[10218] = 8'h16 ;
            rom[10219] = 8'hf6 ;
            rom[10220] = 8'hfc ;
            rom[10221] = 8'h08 ;
            rom[10222] = 8'h03 ;
            rom[10223] = 8'h06 ;
            rom[10224] = 8'he9 ;
            rom[10225] = 8'h06 ;
            rom[10226] = 8'hfe ;
            rom[10227] = 8'h1b ;
            rom[10228] = 8'hd2 ;
            rom[10229] = 8'hf0 ;
            rom[10230] = 8'h14 ;
            rom[10231] = 8'hf9 ;
            rom[10232] = 8'hf1 ;
            rom[10233] = 8'h09 ;
            rom[10234] = 8'h22 ;
            rom[10235] = 8'hec ;
            rom[10236] = 8'hf3 ;
            rom[10237] = 8'h00 ;
            rom[10238] = 8'h1c ;
            rom[10239] = 8'hff ;
            rom[10240] = 8'h20 ;
            rom[10241] = 8'h13 ;
            rom[10242] = 8'hee ;
            rom[10243] = 8'hf6 ;
            rom[10244] = 8'h08 ;
            rom[10245] = 8'h03 ;
            rom[10246] = 8'hff ;
            rom[10247] = 8'hb8 ;
            rom[10248] = 8'hfd ;
            rom[10249] = 8'h08 ;
            rom[10250] = 8'hff ;
            rom[10251] = 8'hd8 ;
            rom[10252] = 8'hd7 ;
            rom[10253] = 8'hf1 ;
            rom[10254] = 8'h1a ;
            rom[10255] = 8'heb ;
            rom[10256] = 8'h13 ;
            rom[10257] = 8'hf2 ;
            rom[10258] = 8'h01 ;
            rom[10259] = 8'hf8 ;
            rom[10260] = 8'he7 ;
            rom[10261] = 8'h04 ;
            rom[10262] = 8'hf7 ;
            rom[10263] = 8'hfc ;
            rom[10264] = 8'hef ;
            rom[10265] = 8'h14 ;
            rom[10266] = 8'h13 ;
            rom[10267] = 8'h05 ;
            rom[10268] = 8'h05 ;
            rom[10269] = 8'hfe ;
            rom[10270] = 8'he0 ;
            rom[10271] = 8'hea ;
            rom[10272] = 8'hf4 ;
            rom[10273] = 8'he6 ;
            rom[10274] = 8'hf0 ;
            rom[10275] = 8'hf8 ;
            rom[10276] = 8'h12 ;
            rom[10277] = 8'h1a ;
            rom[10278] = 8'h09 ;
            rom[10279] = 8'hcd ;
            rom[10280] = 8'hea ;
            rom[10281] = 8'hf8 ;
            rom[10282] = 8'hfc ;
            rom[10283] = 8'h0b ;
            rom[10284] = 8'h12 ;
            rom[10285] = 8'hdd ;
            rom[10286] = 8'hfb ;
            rom[10287] = 8'hde ;
            rom[10288] = 8'hf8 ;
            rom[10289] = 8'h07 ;
            rom[10290] = 8'h0d ;
            rom[10291] = 8'hec ;
            rom[10292] = 8'hef ;
            rom[10293] = 8'hfc ;
            rom[10294] = 8'h07 ;
            rom[10295] = 8'he2 ;
            rom[10296] = 8'he7 ;
            rom[10297] = 8'h00 ;
            rom[10298] = 8'hf9 ;
            rom[10299] = 8'he0 ;
            rom[10300] = 8'hf5 ;
            rom[10301] = 8'h07 ;
            rom[10302] = 8'he3 ;
            rom[10303] = 8'hf4 ;
            rom[10304] = 8'he6 ;
            rom[10305] = 8'hd9 ;
            rom[10306] = 8'hee ;
            rom[10307] = 8'hdd ;
            rom[10308] = 8'h2b ;
            rom[10309] = 8'h10 ;
            rom[10310] = 8'h05 ;
            rom[10311] = 8'hfb ;
            rom[10312] = 8'h19 ;
            rom[10313] = 8'h16 ;
            rom[10314] = 8'h0a ;
            rom[10315] = 8'hbf ;
            rom[10316] = 8'h01 ;
            rom[10317] = 8'h16 ;
            rom[10318] = 8'he4 ;
            rom[10319] = 8'hf0 ;
            rom[10320] = 8'h29 ;
            rom[10321] = 8'h15 ;
            rom[10322] = 8'h07 ;
            rom[10323] = 8'h03 ;
            rom[10324] = 8'he5 ;
            rom[10325] = 8'he1 ;
            rom[10326] = 8'h08 ;
            rom[10327] = 8'h0c ;
            rom[10328] = 8'hef ;
            rom[10329] = 8'h05 ;
            rom[10330] = 8'hfa ;
            rom[10331] = 8'hfa ;
            rom[10332] = 8'h04 ;
            rom[10333] = 8'h02 ;
            rom[10334] = 8'h08 ;
            rom[10335] = 8'heb ;
            rom[10336] = 8'hfd ;
            rom[10337] = 8'hef ;
            rom[10338] = 8'h08 ;
            rom[10339] = 8'h04 ;
            rom[10340] = 8'hd2 ;
            rom[10341] = 8'h14 ;
            rom[10342] = 8'hdd ;
            rom[10343] = 8'hf8 ;
            rom[10344] = 8'h00 ;
            rom[10345] = 8'hff ;
            rom[10346] = 8'h0b ;
            rom[10347] = 8'h05 ;
            rom[10348] = 8'h02 ;
            rom[10349] = 8'hd5 ;
            rom[10350] = 8'he8 ;
            rom[10351] = 8'h07 ;
            rom[10352] = 8'hdd ;
            rom[10353] = 8'h01 ;
            rom[10354] = 8'hf8 ;
            rom[10355] = 8'h05 ;
            rom[10356] = 8'hdb ;
            rom[10357] = 8'hf3 ;
            rom[10358] = 8'hfb ;
            rom[10359] = 8'hf9 ;
            rom[10360] = 8'h02 ;
            rom[10361] = 8'hf2 ;
            rom[10362] = 8'he4 ;
            rom[10363] = 8'h00 ;
            rom[10364] = 8'h15 ;
            rom[10365] = 8'heb ;
            rom[10366] = 8'hea ;
            rom[10367] = 8'h0e ;
            rom[10368] = 8'hf8 ;
            rom[10369] = 8'hea ;
            rom[10370] = 8'h0c ;
            rom[10371] = 8'h10 ;
            rom[10372] = 8'h00 ;
            rom[10373] = 8'he1 ;
            rom[10374] = 8'hcf ;
            rom[10375] = 8'he7 ;
            rom[10376] = 8'h30 ;
            rom[10377] = 8'he9 ;
            rom[10378] = 8'h1b ;
            rom[10379] = 8'h21 ;
            rom[10380] = 8'h1c ;
            rom[10381] = 8'hdc ;
            rom[10382] = 8'hf6 ;
            rom[10383] = 8'hee ;
            rom[10384] = 8'hf2 ;
            rom[10385] = 8'h0b ;
            rom[10386] = 8'hc4 ;
            rom[10387] = 8'h18 ;
            rom[10388] = 8'hff ;
            rom[10389] = 8'hfd ;
            rom[10390] = 8'hea ;
            rom[10391] = 8'hde ;
            rom[10392] = 8'h09 ;
            rom[10393] = 8'h06 ;
            rom[10394] = 8'hdf ;
            rom[10395] = 8'h18 ;
            rom[10396] = 8'hec ;
            rom[10397] = 8'h0c ;
            rom[10398] = 8'hf5 ;
            rom[10399] = 8'hee ;
            rom[10400] = 8'hf8 ;
            rom[10401] = 8'hfd ;
            rom[10402] = 8'h0a ;
            rom[10403] = 8'hf8 ;
            rom[10404] = 8'h13 ;
            rom[10405] = 8'hee ;
            rom[10406] = 8'hfc ;
            rom[10407] = 8'he1 ;
            rom[10408] = 8'hf1 ;
            rom[10409] = 8'hf5 ;
            rom[10410] = 8'hf2 ;
            rom[10411] = 8'hec ;
            rom[10412] = 8'hf8 ;
            rom[10413] = 8'hf4 ;
            rom[10414] = 8'hf2 ;
            rom[10415] = 8'hf5 ;
            rom[10416] = 8'he9 ;
            rom[10417] = 8'hed ;
            rom[10418] = 8'hfe ;
            rom[10419] = 8'h09 ;
            rom[10420] = 8'he7 ;
            rom[10421] = 8'h15 ;
            rom[10422] = 8'h00 ;
            rom[10423] = 8'hf2 ;
            rom[10424] = 8'h01 ;
            rom[10425] = 8'hdd ;
            rom[10426] = 8'hfe ;
            rom[10427] = 8'he5 ;
            rom[10428] = 8'hfa ;
            rom[10429] = 8'hff ;
            rom[10430] = 8'h1c ;
            rom[10431] = 8'hf2 ;
            rom[10432] = 8'h0f ;
            rom[10433] = 8'h12 ;
            rom[10434] = 8'h04 ;
            rom[10435] = 8'h0b ;
            rom[10436] = 8'h00 ;
            rom[10437] = 8'hbc ;
            rom[10438] = 8'hdd ;
            rom[10439] = 8'he9 ;
            rom[10440] = 8'h21 ;
            rom[10441] = 8'he7 ;
            rom[10442] = 8'h16 ;
            rom[10443] = 8'h04 ;
            rom[10444] = 8'he3 ;
            rom[10445] = 8'he9 ;
            rom[10446] = 8'h1e ;
            rom[10447] = 8'h00 ;
            rom[10448] = 8'he3 ;
            rom[10449] = 8'h1e ;
            rom[10450] = 8'h0a ;
            rom[10451] = 8'he6 ;
            rom[10452] = 8'h07 ;
            rom[10453] = 8'he9 ;
            rom[10454] = 8'hec ;
            rom[10455] = 8'hc6 ;
            rom[10456] = 8'h10 ;
            rom[10457] = 8'hf8 ;
            rom[10458] = 8'h0f ;
            rom[10459] = 8'hf7 ;
            rom[10460] = 8'h0b ;
            rom[10461] = 8'h0e ;
            rom[10462] = 8'hf9 ;
            rom[10463] = 8'he5 ;
            rom[10464] = 8'h02 ;
            rom[10465] = 8'h1d ;
            rom[10466] = 8'h00 ;
            rom[10467] = 8'h00 ;
            rom[10468] = 8'hf5 ;
            rom[10469] = 8'hfd ;
            rom[10470] = 8'h18 ;
            rom[10471] = 8'hdc ;
            rom[10472] = 8'hc8 ;
            rom[10473] = 8'h00 ;
            rom[10474] = 8'he7 ;
            rom[10475] = 8'hed ;
            rom[10476] = 8'h09 ;
            rom[10477] = 8'hfb ;
            rom[10478] = 8'h25 ;
            rom[10479] = 8'hea ;
            rom[10480] = 8'h05 ;
            rom[10481] = 8'h01 ;
            rom[10482] = 8'hf6 ;
            rom[10483] = 8'h07 ;
            rom[10484] = 8'h06 ;
            rom[10485] = 8'hf6 ;
            rom[10486] = 8'h1d ;
            rom[10487] = 8'he7 ;
            rom[10488] = 8'h28 ;
            rom[10489] = 8'he8 ;
            rom[10490] = 8'he4 ;
            rom[10491] = 8'h06 ;
            rom[10492] = 8'hfe ;
            rom[10493] = 8'h10 ;
            rom[10494] = 8'h02 ;
            rom[10495] = 8'h04 ;
            rom[10496] = 8'h24 ;
            rom[10497] = 8'h0a ;
            rom[10498] = 8'he9 ;
            rom[10499] = 8'hee ;
            rom[10500] = 8'hf1 ;
            rom[10501] = 8'h03 ;
            rom[10502] = 8'h13 ;
            rom[10503] = 8'h30 ;
            rom[10504] = 8'h04 ;
            rom[10505] = 8'h1a ;
            rom[10506] = 8'hdb ;
            rom[10507] = 8'hef ;
            rom[10508] = 8'he6 ;
            rom[10509] = 8'h05 ;
            rom[10510] = 8'h03 ;
            rom[10511] = 8'hf3 ;
            rom[10512] = 8'hfb ;
            rom[10513] = 8'h13 ;
            rom[10514] = 8'h01 ;
            rom[10515] = 8'h0f ;
            rom[10516] = 8'hf0 ;
            rom[10517] = 8'h01 ;
            rom[10518] = 8'hf7 ;
            rom[10519] = 8'h1a ;
            rom[10520] = 8'hfc ;
            rom[10521] = 8'h06 ;
            rom[10522] = 8'hff ;
            rom[10523] = 8'h14 ;
            rom[10524] = 8'hf7 ;
            rom[10525] = 8'h06 ;
            rom[10526] = 8'h0c ;
            rom[10527] = 8'hf1 ;
            rom[10528] = 8'he9 ;
            rom[10529] = 8'hf3 ;
            rom[10530] = 8'heb ;
            rom[10531] = 8'h13 ;
            rom[10532] = 8'h14 ;
            rom[10533] = 8'h0a ;
            rom[10534] = 8'hcb ;
            rom[10535] = 8'hea ;
            rom[10536] = 8'h07 ;
            rom[10537] = 8'hfd ;
            rom[10538] = 8'hdf ;
            rom[10539] = 8'he8 ;
            rom[10540] = 8'hdf ;
            rom[10541] = 8'he6 ;
            rom[10542] = 8'he2 ;
            rom[10543] = 8'h03 ;
            rom[10544] = 8'he9 ;
            rom[10545] = 8'h13 ;
            rom[10546] = 8'hef ;
            rom[10547] = 8'h06 ;
            rom[10548] = 8'h06 ;
            rom[10549] = 8'hfb ;
            rom[10550] = 8'hf8 ;
            rom[10551] = 8'h03 ;
            rom[10552] = 8'h20 ;
            rom[10553] = 8'hf7 ;
            rom[10554] = 8'h04 ;
            rom[10555] = 8'h0b ;
            rom[10556] = 8'hfa ;
            rom[10557] = 8'h06 ;
            rom[10558] = 8'hed ;
            rom[10559] = 8'hfe ;
            rom[10560] = 8'h2e ;
            rom[10561] = 8'he4 ;
            rom[10562] = 8'h11 ;
            rom[10563] = 8'h03 ;
            rom[10564] = 8'hd8 ;
            rom[10565] = 8'hee ;
            rom[10566] = 8'h0a ;
            rom[10567] = 8'hff ;
            rom[10568] = 8'h00 ;
            rom[10569] = 8'hf6 ;
            rom[10570] = 8'h1a ;
            rom[10571] = 8'h21 ;
            rom[10572] = 8'he1 ;
            rom[10573] = 8'hdb ;
            rom[10574] = 8'hee ;
            rom[10575] = 8'h1f ;
            rom[10576] = 8'hdb ;
            rom[10577] = 8'h09 ;
            rom[10578] = 8'he9 ;
            rom[10579] = 8'he2 ;
            rom[10580] = 8'he7 ;
            rom[10581] = 8'h15 ;
            rom[10582] = 8'h05 ;
            rom[10583] = 8'h28 ;
            rom[10584] = 8'hec ;
            rom[10585] = 8'hea ;
            rom[10586] = 8'hf3 ;
            rom[10587] = 8'hf0 ;
            rom[10588] = 8'he7 ;
            rom[10589] = 8'he1 ;
            rom[10590] = 8'hc6 ;
            rom[10591] = 8'hfb ;
            rom[10592] = 8'hf5 ;
            rom[10593] = 8'h2c ;
            rom[10594] = 8'hd2 ;
            rom[10595] = 8'he5 ;
            rom[10596] = 8'hef ;
            rom[10597] = 8'h01 ;
            rom[10598] = 8'h0a ;
            rom[10599] = 8'h0d ;
            rom[10600] = 8'hc7 ;
            rom[10601] = 8'h0c ;
            rom[10602] = 8'h0c ;
            rom[10603] = 8'hcb ;
            rom[10604] = 8'hf6 ;
            rom[10605] = 8'hfd ;
            rom[10606] = 8'h0f ;
            rom[10607] = 8'h06 ;
            rom[10608] = 8'h21 ;
            rom[10609] = 8'hd3 ;
            rom[10610] = 8'hf7 ;
            rom[10611] = 8'he4 ;
            rom[10612] = 8'h09 ;
            rom[10613] = 8'hf7 ;
            rom[10614] = 8'hf4 ;
            rom[10615] = 8'heb ;
            rom[10616] = 8'hf1 ;
            rom[10617] = 8'h15 ;
            rom[10618] = 8'h00 ;
            rom[10619] = 8'he9 ;
            rom[10620] = 8'h03 ;
            rom[10621] = 8'h10 ;
            rom[10622] = 8'h03 ;
            rom[10623] = 8'hd4 ;
            rom[10624] = 8'hec ;
            rom[10625] = 8'h06 ;
            rom[10626] = 8'hf5 ;
            rom[10627] = 8'h16 ;
            rom[10628] = 8'hde ;
            rom[10629] = 8'hde ;
            rom[10630] = 8'h16 ;
            rom[10631] = 8'h05 ;
            rom[10632] = 8'h19 ;
            rom[10633] = 8'h08 ;
            rom[10634] = 8'h00 ;
            rom[10635] = 8'h00 ;
            rom[10636] = 8'h05 ;
            rom[10637] = 8'hf8 ;
            rom[10638] = 8'he3 ;
            rom[10639] = 8'h0a ;
            rom[10640] = 8'h01 ;
            rom[10641] = 8'h1b ;
            rom[10642] = 8'hd5 ;
            rom[10643] = 8'h08 ;
            rom[10644] = 8'h07 ;
            rom[10645] = 8'hfa ;
            rom[10646] = 8'hef ;
            rom[10647] = 8'hdb ;
            rom[10648] = 8'hf6 ;
            rom[10649] = 8'h14 ;
            rom[10650] = 8'hfe ;
            rom[10651] = 8'h04 ;
            rom[10652] = 8'hc7 ;
            rom[10653] = 8'h1d ;
            rom[10654] = 8'h04 ;
            rom[10655] = 8'hf8 ;
            rom[10656] = 8'h10 ;
            rom[10657] = 8'h06 ;
            rom[10658] = 8'h09 ;
            rom[10659] = 8'hcb ;
            rom[10660] = 8'hef ;
            rom[10661] = 8'hf3 ;
            rom[10662] = 8'hec ;
            rom[10663] = 8'h0c ;
            rom[10664] = 8'h1a ;
            rom[10665] = 8'h13 ;
            rom[10666] = 8'h28 ;
            rom[10667] = 8'h08 ;
            rom[10668] = 8'hf7 ;
            rom[10669] = 8'hbb ;
            rom[10670] = 8'h17 ;
            rom[10671] = 8'hff ;
            rom[10672] = 8'hfc ;
            rom[10673] = 8'h02 ;
            rom[10674] = 8'hd6 ;
            rom[10675] = 8'h15 ;
            rom[10676] = 8'hfd ;
            rom[10677] = 8'hef ;
            rom[10678] = 8'h03 ;
            rom[10679] = 8'hf2 ;
            rom[10680] = 8'he0 ;
            rom[10681] = 8'hf4 ;
            rom[10682] = 8'hb7 ;
            rom[10683] = 8'h04 ;
            rom[10684] = 8'hee ;
            rom[10685] = 8'h02 ;
            rom[10686] = 8'hf5 ;
            rom[10687] = 8'hd6 ;
            rom[10688] = 8'h18 ;
            rom[10689] = 8'hed ;
            rom[10690] = 8'hf9 ;
            rom[10691] = 8'hf0 ;
            rom[10692] = 8'hed ;
            rom[10693] = 8'hdf ;
            rom[10694] = 8'hf8 ;
            rom[10695] = 8'h1a ;
            rom[10696] = 8'h24 ;
            rom[10697] = 8'h12 ;
            rom[10698] = 8'hf4 ;
            rom[10699] = 8'hf6 ;
            rom[10700] = 8'hf5 ;
            rom[10701] = 8'he9 ;
            rom[10702] = 8'h15 ;
            rom[10703] = 8'he3 ;
            rom[10704] = 8'h01 ;
            rom[10705] = 8'h14 ;
            rom[10706] = 8'hf0 ;
            rom[10707] = 8'h02 ;
            rom[10708] = 8'h0b ;
            rom[10709] = 8'hfe ;
            rom[10710] = 8'h02 ;
            rom[10711] = 8'h03 ;
            rom[10712] = 8'he3 ;
            rom[10713] = 8'h11 ;
            rom[10714] = 8'h01 ;
            rom[10715] = 8'hff ;
            rom[10716] = 8'he7 ;
            rom[10717] = 8'h18 ;
            rom[10718] = 8'hef ;
            rom[10719] = 8'hf4 ;
            rom[10720] = 8'h17 ;
            rom[10721] = 8'he8 ;
            rom[10722] = 8'hfc ;
            rom[10723] = 8'hfd ;
            rom[10724] = 8'h12 ;
            rom[10725] = 8'hed ;
            rom[10726] = 8'h07 ;
            rom[10727] = 8'h10 ;
            rom[10728] = 8'hef ;
            rom[10729] = 8'h01 ;
            rom[10730] = 8'hec ;
            rom[10731] = 8'h07 ;
            rom[10732] = 8'hf7 ;
            rom[10733] = 8'h03 ;
            rom[10734] = 8'h02 ;
            rom[10735] = 8'hf7 ;
            rom[10736] = 8'hfc ;
            rom[10737] = 8'he4 ;
            rom[10738] = 8'hfc ;
            rom[10739] = 8'he4 ;
            rom[10740] = 8'h00 ;
            rom[10741] = 8'h06 ;
            rom[10742] = 8'he9 ;
            rom[10743] = 8'he1 ;
            rom[10744] = 8'h01 ;
            rom[10745] = 8'h00 ;
            rom[10746] = 8'he9 ;
            rom[10747] = 8'h01 ;
            rom[10748] = 8'h08 ;
            rom[10749] = 8'hd9 ;
            rom[10750] = 8'h25 ;
            rom[10751] = 8'hd8 ;
            rom[10752] = 8'h07 ;
            rom[10753] = 8'he8 ;
            rom[10754] = 8'hf7 ;
            rom[10755] = 8'hc1 ;
            rom[10756] = 8'hd9 ;
            rom[10757] = 8'h01 ;
            rom[10758] = 8'h01 ;
            rom[10759] = 8'hf9 ;
            rom[10760] = 8'h12 ;
            rom[10761] = 8'h06 ;
            rom[10762] = 8'hf1 ;
            rom[10763] = 8'he5 ;
            rom[10764] = 8'h09 ;
            rom[10765] = 8'h0e ;
            rom[10766] = 8'h0a ;
            rom[10767] = 8'h0b ;
            rom[10768] = 8'h01 ;
            rom[10769] = 8'h0f ;
            rom[10770] = 8'h18 ;
            rom[10771] = 8'hf3 ;
            rom[10772] = 8'hc1 ;
            rom[10773] = 8'hfa ;
            rom[10774] = 8'h07 ;
            rom[10775] = 8'h0d ;
            rom[10776] = 8'hf0 ;
            rom[10777] = 8'h01 ;
            rom[10778] = 8'h09 ;
            rom[10779] = 8'hfb ;
            rom[10780] = 8'h04 ;
            rom[10781] = 8'he2 ;
            rom[10782] = 8'hfb ;
            rom[10783] = 8'hd8 ;
            rom[10784] = 8'hf8 ;
            rom[10785] = 8'hf7 ;
            rom[10786] = 8'h07 ;
            rom[10787] = 8'h04 ;
            rom[10788] = 8'hf3 ;
            rom[10789] = 8'h1c ;
            rom[10790] = 8'h09 ;
            rom[10791] = 8'hf5 ;
            rom[10792] = 8'he9 ;
            rom[10793] = 8'h17 ;
            rom[10794] = 8'h18 ;
            rom[10795] = 8'he9 ;
            rom[10796] = 8'h04 ;
            rom[10797] = 8'hf7 ;
            rom[10798] = 8'h10 ;
            rom[10799] = 8'h0e ;
            rom[10800] = 8'h08 ;
            rom[10801] = 8'hf4 ;
            rom[10802] = 8'hbc ;
            rom[10803] = 8'h21 ;
            rom[10804] = 8'h0a ;
            rom[10805] = 8'hfe ;
            rom[10806] = 8'hf6 ;
            rom[10807] = 8'hdd ;
            rom[10808] = 8'h02 ;
            rom[10809] = 8'hfd ;
            rom[10810] = 8'hff ;
            rom[10811] = 8'h0d ;
            rom[10812] = 8'h03 ;
            rom[10813] = 8'hf4 ;
            rom[10814] = 8'h01 ;
            rom[10815] = 8'h1c ;
            rom[10816] = 8'h13 ;
            rom[10817] = 8'hf7 ;
            rom[10818] = 8'hec ;
            rom[10819] = 8'he6 ;
            rom[10820] = 8'hf8 ;
            rom[10821] = 8'h11 ;
            rom[10822] = 8'h06 ;
            rom[10823] = 8'hf9 ;
            rom[10824] = 8'h19 ;
            rom[10825] = 8'h01 ;
            rom[10826] = 8'h0c ;
            rom[10827] = 8'he9 ;
            rom[10828] = 8'h13 ;
            rom[10829] = 8'h16 ;
            rom[10830] = 8'h0f ;
            rom[10831] = 8'hec ;
            rom[10832] = 8'hf3 ;
            rom[10833] = 8'h02 ;
            rom[10834] = 8'h05 ;
            rom[10835] = 8'h01 ;
            rom[10836] = 8'hf7 ;
            rom[10837] = 8'hf3 ;
            rom[10838] = 8'h1f ;
            rom[10839] = 8'hfb ;
            rom[10840] = 8'h07 ;
            rom[10841] = 8'hea ;
            rom[10842] = 8'hfe ;
            rom[10843] = 8'hef ;
            rom[10844] = 8'hfc ;
            rom[10845] = 8'hf3 ;
            rom[10846] = 8'h1c ;
            rom[10847] = 8'hec ;
            rom[10848] = 8'hf3 ;
            rom[10849] = 8'h0d ;
            rom[10850] = 8'h18 ;
            rom[10851] = 8'hfb ;
            rom[10852] = 8'hee ;
            rom[10853] = 8'h25 ;
            rom[10854] = 8'hee ;
            rom[10855] = 8'hf7 ;
            rom[10856] = 8'h17 ;
            rom[10857] = 8'h13 ;
            rom[10858] = 8'h2b ;
            rom[10859] = 8'h0a ;
            rom[10860] = 8'h1b ;
            rom[10861] = 8'he6 ;
            rom[10862] = 8'h06 ;
            rom[10863] = 8'h08 ;
            rom[10864] = 8'hdf ;
            rom[10865] = 8'h01 ;
            rom[10866] = 8'hab ;
            rom[10867] = 8'h11 ;
            rom[10868] = 8'he6 ;
            rom[10869] = 8'hf4 ;
            rom[10870] = 8'h0c ;
            rom[10871] = 8'hd1 ;
            rom[10872] = 8'h08 ;
            rom[10873] = 8'hf6 ;
            rom[10874] = 8'he0 ;
            rom[10875] = 8'h08 ;
            rom[10876] = 8'h11 ;
            rom[10877] = 8'hf1 ;
            rom[10878] = 8'h01 ;
            rom[10879] = 8'h2c ;
            rom[10880] = 8'hf1 ;
            rom[10881] = 8'hcc ;
            rom[10882] = 8'h15 ;
            rom[10883] = 8'hfc ;
            rom[10884] = 8'hfc ;
            rom[10885] = 8'h0d ;
            rom[10886] = 8'h15 ;
            rom[10887] = 8'hd0 ;
            rom[10888] = 8'h10 ;
            rom[10889] = 8'hf3 ;
            rom[10890] = 8'h04 ;
            rom[10891] = 8'h04 ;
            rom[10892] = 8'hf5 ;
            rom[10893] = 8'h02 ;
            rom[10894] = 8'h11 ;
            rom[10895] = 8'h0a ;
            rom[10896] = 8'hf0 ;
            rom[10897] = 8'h05 ;
            rom[10898] = 8'h07 ;
            rom[10899] = 8'h11 ;
            rom[10900] = 8'h11 ;
            rom[10901] = 8'h1a ;
            rom[10902] = 8'h0d ;
            rom[10903] = 8'hf1 ;
            rom[10904] = 8'hfb ;
            rom[10905] = 8'hf9 ;
            rom[10906] = 8'h12 ;
            rom[10907] = 8'hd2 ;
            rom[10908] = 8'hec ;
            rom[10909] = 8'hfd ;
            rom[10910] = 8'h05 ;
            rom[10911] = 8'he2 ;
            rom[10912] = 8'hfa ;
            rom[10913] = 8'h05 ;
            rom[10914] = 8'h05 ;
            rom[10915] = 8'hfb ;
            rom[10916] = 8'h00 ;
            rom[10917] = 8'h0c ;
            rom[10918] = 8'h1c ;
            rom[10919] = 8'h0d ;
            rom[10920] = 8'hdd ;
            rom[10921] = 8'h13 ;
            rom[10922] = 8'h0c ;
            rom[10923] = 8'hfb ;
            rom[10924] = 8'h20 ;
            rom[10925] = 8'hfd ;
            rom[10926] = 8'h17 ;
            rom[10927] = 8'h20 ;
            rom[10928] = 8'hd8 ;
            rom[10929] = 8'hfb ;
            rom[10930] = 8'h00 ;
            rom[10931] = 8'hec ;
            rom[10932] = 8'h18 ;
            rom[10933] = 8'hfb ;
            rom[10934] = 8'hd7 ;
            rom[10935] = 8'hef ;
            rom[10936] = 8'hf6 ;
            rom[10937] = 8'h0a ;
            rom[10938] = 8'hf0 ;
            rom[10939] = 8'hfd ;
            rom[10940] = 8'h0a ;
            rom[10941] = 8'h18 ;
            rom[10942] = 8'h08 ;
            rom[10943] = 8'hec ;
            rom[10944] = 8'hfa ;
            rom[10945] = 8'h1d ;
            rom[10946] = 8'h17 ;
            rom[10947] = 8'he5 ;
            rom[10948] = 8'he0 ;
            rom[10949] = 8'h08 ;
            rom[10950] = 8'h08 ;
            rom[10951] = 8'hf5 ;
            rom[10952] = 8'h14 ;
            rom[10953] = 8'h12 ;
            rom[10954] = 8'hf1 ;
            rom[10955] = 8'h15 ;
            rom[10956] = 8'h0f ;
            rom[10957] = 8'hea ;
            rom[10958] = 8'h20 ;
            rom[10959] = 8'h08 ;
            rom[10960] = 8'h05 ;
            rom[10961] = 8'hd9 ;
            rom[10962] = 8'h00 ;
            rom[10963] = 8'hf7 ;
            rom[10964] = 8'hfb ;
            rom[10965] = 8'h09 ;
            rom[10966] = 8'hff ;
            rom[10967] = 8'hff ;
            rom[10968] = 8'h06 ;
            rom[10969] = 8'he3 ;
            rom[10970] = 8'h16 ;
            rom[10971] = 8'h0f ;
            rom[10972] = 8'h1b ;
            rom[10973] = 8'hf0 ;
            rom[10974] = 8'h2a ;
            rom[10975] = 8'hfe ;
            rom[10976] = 8'h03 ;
            rom[10977] = 8'hf5 ;
            rom[10978] = 8'h1a ;
            rom[10979] = 8'hee ;
            rom[10980] = 8'hdd ;
            rom[10981] = 8'h16 ;
            rom[10982] = 8'hee ;
            rom[10983] = 8'h03 ;
            rom[10984] = 8'hd9 ;
            rom[10985] = 8'h00 ;
            rom[10986] = 8'he6 ;
            rom[10987] = 8'he1 ;
            rom[10988] = 8'hee ;
            rom[10989] = 8'hef ;
            rom[10990] = 8'he0 ;
            rom[10991] = 8'h19 ;
            rom[10992] = 8'hea ;
            rom[10993] = 8'hdd ;
            rom[10994] = 8'h14 ;
            rom[10995] = 8'hfc ;
            rom[10996] = 8'h14 ;
            rom[10997] = 8'hfc ;
            rom[10998] = 8'h0f ;
            rom[10999] = 8'h1d ;
            rom[11000] = 8'h11 ;
            rom[11001] = 8'h15 ;
            rom[11002] = 8'he2 ;
            rom[11003] = 8'he5 ;
            rom[11004] = 8'hfe ;
            rom[11005] = 8'h0d ;
            rom[11006] = 8'h0a ;
            rom[11007] = 8'h08 ;
            rom[11008] = 8'hf3 ;
            rom[11009] = 8'h0e ;
            rom[11010] = 8'h07 ;
            rom[11011] = 8'hf2 ;
            rom[11012] = 8'hed ;
            rom[11013] = 8'h03 ;
            rom[11014] = 8'hfe ;
            rom[11015] = 8'hfd ;
            rom[11016] = 8'h30 ;
            rom[11017] = 8'h14 ;
            rom[11018] = 8'h0d ;
            rom[11019] = 8'heb ;
            rom[11020] = 8'h07 ;
            rom[11021] = 8'h00 ;
            rom[11022] = 8'he9 ;
            rom[11023] = 8'h11 ;
            rom[11024] = 8'hfd ;
            rom[11025] = 8'h0a ;
            rom[11026] = 8'he4 ;
            rom[11027] = 8'h06 ;
            rom[11028] = 8'hef ;
            rom[11029] = 8'h0e ;
            rom[11030] = 8'hfb ;
            rom[11031] = 8'he5 ;
            rom[11032] = 8'hcb ;
            rom[11033] = 8'h05 ;
            rom[11034] = 8'hed ;
            rom[11035] = 8'hfc ;
            rom[11036] = 8'hc8 ;
            rom[11037] = 8'h0b ;
            rom[11038] = 8'h21 ;
            rom[11039] = 8'hfb ;
            rom[11040] = 8'h39 ;
            rom[11041] = 8'hf2 ;
            rom[11042] = 8'h00 ;
            rom[11043] = 8'hfc ;
            rom[11044] = 8'hea ;
            rom[11045] = 8'hf6 ;
            rom[11046] = 8'hca ;
            rom[11047] = 8'h0b ;
            rom[11048] = 8'h13 ;
            rom[11049] = 8'h00 ;
            rom[11050] = 8'h15 ;
            rom[11051] = 8'h17 ;
            rom[11052] = 8'hfb ;
            rom[11053] = 8'hb7 ;
            rom[11054] = 8'h04 ;
            rom[11055] = 8'h12 ;
            rom[11056] = 8'he3 ;
            rom[11057] = 8'hec ;
            rom[11058] = 8'hec ;
            rom[11059] = 8'h01 ;
            rom[11060] = 8'hf7 ;
            rom[11061] = 8'he6 ;
            rom[11062] = 8'hff ;
            rom[11063] = 8'heb ;
            rom[11064] = 8'h12 ;
            rom[11065] = 8'he7 ;
            rom[11066] = 8'hcb ;
            rom[11067] = 8'hfe ;
            rom[11068] = 8'h0a ;
            rom[11069] = 8'he9 ;
            rom[11070] = 8'h06 ;
            rom[11071] = 8'hde ;
            rom[11072] = 8'hfa ;
            rom[11073] = 8'h13 ;
            rom[11074] = 8'hef ;
            rom[11075] = 8'he3 ;
            rom[11076] = 8'hd9 ;
            rom[11077] = 8'h0e ;
            rom[11078] = 8'h0d ;
            rom[11079] = 8'h0d ;
            rom[11080] = 8'h09 ;
            rom[11081] = 8'h0d ;
            rom[11082] = 8'hf0 ;
            rom[11083] = 8'hc3 ;
            rom[11084] = 8'hce ;
            rom[11085] = 8'hf1 ;
            rom[11086] = 8'h12 ;
            rom[11087] = 8'h0f ;
            rom[11088] = 8'h04 ;
            rom[11089] = 8'hfa ;
            rom[11090] = 8'h0a ;
            rom[11091] = 8'hcf ;
            rom[11092] = 8'he1 ;
            rom[11093] = 8'h04 ;
            rom[11094] = 8'h08 ;
            rom[11095] = 8'h15 ;
            rom[11096] = 8'h0b ;
            rom[11097] = 8'hff ;
            rom[11098] = 8'h00 ;
            rom[11099] = 8'h07 ;
            rom[11100] = 8'hfa ;
            rom[11101] = 8'hfb ;
            rom[11102] = 8'h03 ;
            rom[11103] = 8'hfa ;
            rom[11104] = 8'hdc ;
            rom[11105] = 8'hec ;
            rom[11106] = 8'hf0 ;
            rom[11107] = 8'h1c ;
            rom[11108] = 8'h10 ;
            rom[11109] = 8'h0f ;
            rom[11110] = 8'hf8 ;
            rom[11111] = 8'he9 ;
            rom[11112] = 8'he3 ;
            rom[11113] = 8'h16 ;
            rom[11114] = 8'hef ;
            rom[11115] = 8'hf4 ;
            rom[11116] = 8'hf1 ;
            rom[11117] = 8'hee ;
            rom[11118] = 8'hfa ;
            rom[11119] = 8'he7 ;
            rom[11120] = 8'h1a ;
            rom[11121] = 8'hf4 ;
            rom[11122] = 8'h14 ;
            rom[11123] = 8'hfc ;
            rom[11124] = 8'hed ;
            rom[11125] = 8'hfd ;
            rom[11126] = 8'hf7 ;
            rom[11127] = 8'hdd ;
            rom[11128] = 8'hf6 ;
            rom[11129] = 8'hff ;
            rom[11130] = 8'h05 ;
            rom[11131] = 8'hf0 ;
            rom[11132] = 8'hf0 ;
            rom[11133] = 8'he7 ;
            rom[11134] = 8'he2 ;
            rom[11135] = 8'he2 ;
            rom[11136] = 8'h1e ;
            rom[11137] = 8'h06 ;
            rom[11138] = 8'hef ;
            rom[11139] = 8'hfd ;
            rom[11140] = 8'hea ;
            rom[11141] = 8'hed ;
            rom[11142] = 8'hff ;
            rom[11143] = 8'he1 ;
            rom[11144] = 8'h1d ;
            rom[11145] = 8'hf5 ;
            rom[11146] = 8'h05 ;
            rom[11147] = 8'h11 ;
            rom[11148] = 8'hf8 ;
            rom[11149] = 8'hfc ;
            rom[11150] = 8'h0b ;
            rom[11151] = 8'hf1 ;
            rom[11152] = 8'h09 ;
            rom[11153] = 8'hfa ;
            rom[11154] = 8'hf5 ;
            rom[11155] = 8'hfc ;
            rom[11156] = 8'h00 ;
            rom[11157] = 8'h0c ;
            rom[11158] = 8'hcd ;
            rom[11159] = 8'hc8 ;
            rom[11160] = 8'h07 ;
            rom[11161] = 8'h0a ;
            rom[11162] = 8'he9 ;
            rom[11163] = 8'h0a ;
            rom[11164] = 8'h0f ;
            rom[11165] = 8'h0b ;
            rom[11166] = 8'h01 ;
            rom[11167] = 8'hed ;
            rom[11168] = 8'h15 ;
            rom[11169] = 8'h36 ;
            rom[11170] = 8'h06 ;
            rom[11171] = 8'h26 ;
            rom[11172] = 8'hf4 ;
            rom[11173] = 8'h19 ;
            rom[11174] = 8'hfb ;
            rom[11175] = 8'hf8 ;
            rom[11176] = 8'h02 ;
            rom[11177] = 8'h0b ;
            rom[11178] = 8'h12 ;
            rom[11179] = 8'h18 ;
            rom[11180] = 8'hf3 ;
            rom[11181] = 8'hc6 ;
            rom[11182] = 8'hff ;
            rom[11183] = 8'he9 ;
            rom[11184] = 8'hf7 ;
            rom[11185] = 8'hfb ;
            rom[11186] = 8'h18 ;
            rom[11187] = 8'h07 ;
            rom[11188] = 8'he7 ;
            rom[11189] = 8'hf2 ;
            rom[11190] = 8'hf5 ;
            rom[11191] = 8'he0 ;
            rom[11192] = 8'h15 ;
            rom[11193] = 8'h1a ;
            rom[11194] = 8'hfc ;
            rom[11195] = 8'hef ;
            rom[11196] = 8'h09 ;
            rom[11197] = 8'hfe ;
            rom[11198] = 8'hfa ;
            rom[11199] = 8'he9 ;
            rom[11200] = 8'h0a ;
            rom[11201] = 8'hfd ;
            rom[11202] = 8'h13 ;
            rom[11203] = 8'h0a ;
            rom[11204] = 8'hed ;
            rom[11205] = 8'h10 ;
            rom[11206] = 8'hfe ;
            rom[11207] = 8'he9 ;
            rom[11208] = 8'h1d ;
            rom[11209] = 8'hfd ;
            rom[11210] = 8'h09 ;
            rom[11211] = 8'hee ;
            rom[11212] = 8'hf2 ;
            rom[11213] = 8'hf6 ;
            rom[11214] = 8'hed ;
            rom[11215] = 8'h02 ;
            rom[11216] = 8'hfb ;
            rom[11217] = 8'hc7 ;
            rom[11218] = 8'hc3 ;
            rom[11219] = 8'he8 ;
            rom[11220] = 8'h08 ;
            rom[11221] = 8'hf8 ;
            rom[11222] = 8'hf3 ;
            rom[11223] = 8'h04 ;
            rom[11224] = 8'h07 ;
            rom[11225] = 8'hfe ;
            rom[11226] = 8'hee ;
            rom[11227] = 8'h15 ;
            rom[11228] = 8'h04 ;
            rom[11229] = 8'h05 ;
            rom[11230] = 8'h29 ;
            rom[11231] = 8'hf5 ;
            rom[11232] = 8'h09 ;
            rom[11233] = 8'h19 ;
            rom[11234] = 8'h02 ;
            rom[11235] = 8'h03 ;
            rom[11236] = 8'h0e ;
            rom[11237] = 8'h1b ;
            rom[11238] = 8'he2 ;
            rom[11239] = 8'h02 ;
            rom[11240] = 8'h22 ;
            rom[11241] = 8'h0a ;
            rom[11242] = 8'hf3 ;
            rom[11243] = 8'h0f ;
            rom[11244] = 8'he3 ;
            rom[11245] = 8'hcb ;
            rom[11246] = 8'hec ;
            rom[11247] = 8'h16 ;
            rom[11248] = 8'hd2 ;
            rom[11249] = 8'hdd ;
            rom[11250] = 8'h14 ;
            rom[11251] = 8'hf0 ;
            rom[11252] = 8'h00 ;
            rom[11253] = 8'h00 ;
            rom[11254] = 8'h01 ;
            rom[11255] = 8'hee ;
            rom[11256] = 8'h11 ;
            rom[11257] = 8'hf4 ;
            rom[11258] = 8'hcc ;
            rom[11259] = 8'hee ;
            rom[11260] = 8'hea ;
            rom[11261] = 8'h07 ;
            rom[11262] = 8'h2b ;
            rom[11263] = 8'h0c ;
            rom[11264] = 8'h0c ;
            rom[11265] = 8'h14 ;
            rom[11266] = 8'hf5 ;
            rom[11267] = 8'h13 ;
            rom[11268] = 8'hf0 ;
            rom[11269] = 8'he4 ;
            rom[11270] = 8'h03 ;
            rom[11271] = 8'hef ;
            rom[11272] = 8'h11 ;
            rom[11273] = 8'h06 ;
            rom[11274] = 8'h05 ;
            rom[11275] = 8'he1 ;
            rom[11276] = 8'h11 ;
            rom[11277] = 8'hda ;
            rom[11278] = 8'hdb ;
            rom[11279] = 8'h17 ;
            rom[11280] = 8'h09 ;
            rom[11281] = 8'h13 ;
            rom[11282] = 8'h06 ;
            rom[11283] = 8'h16 ;
            rom[11284] = 8'hfc ;
            rom[11285] = 8'hfd ;
            rom[11286] = 8'hfc ;
            rom[11287] = 8'he5 ;
            rom[11288] = 8'hf6 ;
            rom[11289] = 8'h08 ;
            rom[11290] = 8'he4 ;
            rom[11291] = 8'hfa ;
            rom[11292] = 8'hb4 ;
            rom[11293] = 8'h12 ;
            rom[11294] = 8'hff ;
            rom[11295] = 8'h0c ;
            rom[11296] = 8'h20 ;
            rom[11297] = 8'h27 ;
            rom[11298] = 8'h07 ;
            rom[11299] = 8'he2 ;
            rom[11300] = 8'hef ;
            rom[11301] = 8'hfc ;
            rom[11302] = 8'h08 ;
            rom[11303] = 8'hef ;
            rom[11304] = 8'h0d ;
            rom[11305] = 8'h14 ;
            rom[11306] = 8'h01 ;
            rom[11307] = 8'h17 ;
            rom[11308] = 8'hf0 ;
            rom[11309] = 8'hd6 ;
            rom[11310] = 8'h22 ;
            rom[11311] = 8'h0a ;
            rom[11312] = 8'h0d ;
            rom[11313] = 8'hfa ;
            rom[11314] = 8'h10 ;
            rom[11315] = 8'hfb ;
            rom[11316] = 8'h00 ;
            rom[11317] = 8'hd1 ;
            rom[11318] = 8'h09 ;
            rom[11319] = 8'hef ;
            rom[11320] = 8'hfb ;
            rom[11321] = 8'heb ;
            rom[11322] = 8'hf7 ;
            rom[11323] = 8'h01 ;
            rom[11324] = 8'hf1 ;
            rom[11325] = 8'h14 ;
            rom[11326] = 8'hfe ;
            rom[11327] = 8'hdd ;
            rom[11328] = 8'he0 ;
            rom[11329] = 8'hef ;
            rom[11330] = 8'hd6 ;
            rom[11331] = 8'hf5 ;
            rom[11332] = 8'h23 ;
            rom[11333] = 8'h02 ;
            rom[11334] = 8'h02 ;
            rom[11335] = 8'h0f ;
            rom[11336] = 8'h05 ;
            rom[11337] = 8'h2c ;
            rom[11338] = 8'he0 ;
            rom[11339] = 8'hf1 ;
            rom[11340] = 8'h04 ;
            rom[11341] = 8'h12 ;
            rom[11342] = 8'hfa ;
            rom[11343] = 8'hed ;
            rom[11344] = 8'h15 ;
            rom[11345] = 8'h13 ;
            rom[11346] = 8'h14 ;
            rom[11347] = 8'hf8 ;
            rom[11348] = 8'h0f ;
            rom[11349] = 8'h03 ;
            rom[11350] = 8'hf5 ;
            rom[11351] = 8'h00 ;
            rom[11352] = 8'hfc ;
            rom[11353] = 8'h03 ;
            rom[11354] = 8'h06 ;
            rom[11355] = 8'he1 ;
            rom[11356] = 8'h06 ;
            rom[11357] = 8'h06 ;
            rom[11358] = 8'hfc ;
            rom[11359] = 8'hfa ;
            rom[11360] = 8'h0f ;
            rom[11361] = 8'he8 ;
            rom[11362] = 8'hfa ;
            rom[11363] = 8'hf7 ;
            rom[11364] = 8'h15 ;
            rom[11365] = 8'h00 ;
            rom[11366] = 8'h01 ;
            rom[11367] = 8'hd8 ;
            rom[11368] = 8'hdd ;
            rom[11369] = 8'hff ;
            rom[11370] = 8'hf5 ;
            rom[11371] = 8'hd4 ;
            rom[11372] = 8'h0c ;
            rom[11373] = 8'hfd ;
            rom[11374] = 8'heb ;
            rom[11375] = 8'hf8 ;
            rom[11376] = 8'hfd ;
            rom[11377] = 8'hfb ;
            rom[11378] = 8'he6 ;
            rom[11379] = 8'h11 ;
            rom[11380] = 8'h1a ;
            rom[11381] = 8'hf6 ;
            rom[11382] = 8'h0b ;
            rom[11383] = 8'hf7 ;
            rom[11384] = 8'hf0 ;
            rom[11385] = 8'h00 ;
            rom[11386] = 8'hfa ;
            rom[11387] = 8'h0d ;
            rom[11388] = 8'h06 ;
            rom[11389] = 8'he6 ;
            rom[11390] = 8'h06 ;
            rom[11391] = 8'h0e ;
            rom[11392] = 8'h0b ;
            rom[11393] = 8'h02 ;
            rom[11394] = 8'hcc ;
            rom[11395] = 8'h00 ;
            rom[11396] = 8'hed ;
            rom[11397] = 8'he8 ;
            rom[11398] = 8'h2e ;
            rom[11399] = 8'h0e ;
            rom[11400] = 8'h13 ;
            rom[11401] = 8'h0d ;
            rom[11402] = 8'h00 ;
            rom[11403] = 8'hfc ;
            rom[11404] = 8'hf8 ;
            rom[11405] = 8'hb9 ;
            rom[11406] = 8'hfb ;
            rom[11407] = 8'h01 ;
            rom[11408] = 8'hf8 ;
            rom[11409] = 8'h15 ;
            rom[11410] = 8'hfa ;
            rom[11411] = 8'h10 ;
            rom[11412] = 8'hfb ;
            rom[11413] = 8'h18 ;
            rom[11414] = 8'h1e ;
            rom[11415] = 8'hf1 ;
            rom[11416] = 8'h05 ;
            rom[11417] = 8'hf9 ;
            rom[11418] = 8'h19 ;
            rom[11419] = 8'h01 ;
            rom[11420] = 8'he9 ;
            rom[11421] = 8'hf8 ;
            rom[11422] = 8'h0c ;
            rom[11423] = 8'hdc ;
            rom[11424] = 8'h19 ;
            rom[11425] = 8'hf9 ;
            rom[11426] = 8'hdc ;
            rom[11427] = 8'h04 ;
            rom[11428] = 8'h02 ;
            rom[11429] = 8'hec ;
            rom[11430] = 8'h00 ;
            rom[11431] = 8'h15 ;
            rom[11432] = 8'h07 ;
            rom[11433] = 8'h15 ;
            rom[11434] = 8'h10 ;
            rom[11435] = 8'h12 ;
            rom[11436] = 8'he7 ;
            rom[11437] = 8'hdf ;
            rom[11438] = 8'h1c ;
            rom[11439] = 8'he4 ;
            rom[11440] = 8'hf3 ;
            rom[11441] = 8'h0b ;
            rom[11442] = 8'hf5 ;
            rom[11443] = 8'h02 ;
            rom[11444] = 8'hf8 ;
            rom[11445] = 8'hd8 ;
            rom[11446] = 8'h0b ;
            rom[11447] = 8'hf6 ;
            rom[11448] = 8'h10 ;
            rom[11449] = 8'he7 ;
            rom[11450] = 8'hfc ;
            rom[11451] = 8'h07 ;
            rom[11452] = 8'h02 ;
            rom[11453] = 8'h24 ;
            rom[11454] = 8'hda ;
            rom[11455] = 8'hc9 ;
            rom[11456] = 8'hf4 ;
            rom[11457] = 8'h35 ;
            rom[11458] = 8'hf7 ;
            rom[11459] = 8'hbd ;
            rom[11460] = 8'hda ;
            rom[11461] = 8'hef ;
            rom[11462] = 8'hf3 ;
            rom[11463] = 8'h01 ;
            rom[11464] = 8'hea ;
            rom[11465] = 8'hf3 ;
            rom[11466] = 8'hba ;
            rom[11467] = 8'hf0 ;
            rom[11468] = 8'he6 ;
            rom[11469] = 8'h00 ;
            rom[11470] = 8'h01 ;
            rom[11471] = 8'h07 ;
            rom[11472] = 8'hf3 ;
            rom[11473] = 8'hff ;
            rom[11474] = 8'h11 ;
            rom[11475] = 8'he2 ;
            rom[11476] = 8'hac ;
            rom[11477] = 8'h15 ;
            rom[11478] = 8'hff ;
            rom[11479] = 8'h15 ;
            rom[11480] = 8'h07 ;
            rom[11481] = 8'h01 ;
            rom[11482] = 8'h05 ;
            rom[11483] = 8'h0d ;
            rom[11484] = 8'hf0 ;
            rom[11485] = 8'h01 ;
            rom[11486] = 8'h0d ;
            rom[11487] = 8'hd9 ;
            rom[11488] = 8'h07 ;
            rom[11489] = 8'hb6 ;
            rom[11490] = 8'hf3 ;
            rom[11491] = 8'h07 ;
            rom[11492] = 8'hfa ;
            rom[11493] = 8'h10 ;
            rom[11494] = 8'hd8 ;
            rom[11495] = 8'he7 ;
            rom[11496] = 8'hf7 ;
            rom[11497] = 8'hf3 ;
            rom[11498] = 8'hf1 ;
            rom[11499] = 8'he9 ;
            rom[11500] = 8'hf7 ;
            rom[11501] = 8'h0d ;
            rom[11502] = 8'hca ;
            rom[11503] = 8'h06 ;
            rom[11504] = 8'h05 ;
            rom[11505] = 8'he9 ;
            rom[11506] = 8'hf3 ;
            rom[11507] = 8'h10 ;
            rom[11508] = 8'h00 ;
            rom[11509] = 8'h0c ;
            rom[11510] = 8'hec ;
            rom[11511] = 8'hfc ;
            rom[11512] = 8'hf2 ;
            rom[11513] = 8'h30 ;
            rom[11514] = 8'hf0 ;
            rom[11515] = 8'hed ;
            rom[11516] = 8'hf9 ;
            rom[11517] = 8'h0b ;
            rom[11518] = 8'h19 ;
            rom[11519] = 8'h17 ;
            rom[11520] = 8'hf4 ;
            rom[11521] = 8'h15 ;
            rom[11522] = 8'hde ;
            rom[11523] = 8'hfc ;
            rom[11524] = 8'hf5 ;
            rom[11525] = 8'hfe ;
            rom[11526] = 8'h05 ;
            rom[11527] = 8'hf8 ;
            rom[11528] = 8'h0a ;
            rom[11529] = 8'h20 ;
            rom[11530] = 8'hfc ;
            rom[11531] = 8'h05 ;
            rom[11532] = 8'h20 ;
            rom[11533] = 8'h08 ;
            rom[11534] = 8'hd6 ;
            rom[11535] = 8'h18 ;
            rom[11536] = 8'h12 ;
            rom[11537] = 8'h17 ;
            rom[11538] = 8'h24 ;
            rom[11539] = 8'h05 ;
            rom[11540] = 8'hd1 ;
            rom[11541] = 8'h04 ;
            rom[11542] = 8'h01 ;
            rom[11543] = 8'hf2 ;
            rom[11544] = 8'hfd ;
            rom[11545] = 8'h10 ;
            rom[11546] = 8'h10 ;
            rom[11547] = 8'he1 ;
            rom[11548] = 8'h0e ;
            rom[11549] = 8'hfb ;
            rom[11550] = 8'hfb ;
            rom[11551] = 8'h02 ;
            rom[11552] = 8'h08 ;
            rom[11553] = 8'h03 ;
            rom[11554] = 8'h0e ;
            rom[11555] = 8'he4 ;
            rom[11556] = 8'hfb ;
            rom[11557] = 8'h08 ;
            rom[11558] = 8'h14 ;
            rom[11559] = 8'hf7 ;
            rom[11560] = 8'h12 ;
            rom[11561] = 8'h17 ;
            rom[11562] = 8'h03 ;
            rom[11563] = 8'h0d ;
            rom[11564] = 8'hfd ;
            rom[11565] = 8'hf4 ;
            rom[11566] = 8'h06 ;
            rom[11567] = 8'hd8 ;
            rom[11568] = 8'h0e ;
            rom[11569] = 8'hf8 ;
            rom[11570] = 8'hc4 ;
            rom[11571] = 8'h20 ;
            rom[11572] = 8'h0d ;
            rom[11573] = 8'hdc ;
            rom[11574] = 8'h02 ;
            rom[11575] = 8'hf4 ;
            rom[11576] = 8'h09 ;
            rom[11577] = 8'hd0 ;
            rom[11578] = 8'h03 ;
            rom[11579] = 8'h09 ;
            rom[11580] = 8'h06 ;
            rom[11581] = 8'h09 ;
            rom[11582] = 8'hd9 ;
            rom[11583] = 8'h06 ;
            rom[11584] = 8'h0a ;
            rom[11585] = 8'he1 ;
            rom[11586] = 8'h1c ;
            rom[11587] = 8'h11 ;
            rom[11588] = 8'hdc ;
            rom[11589] = 8'hcc ;
            rom[11590] = 8'hf0 ;
            rom[11591] = 8'h18 ;
            rom[11592] = 8'h1b ;
            rom[11593] = 8'hdd ;
            rom[11594] = 8'h19 ;
            rom[11595] = 8'h19 ;
            rom[11596] = 8'hfc ;
            rom[11597] = 8'hf1 ;
            rom[11598] = 8'h0d ;
            rom[11599] = 8'h1d ;
            rom[11600] = 8'h02 ;
            rom[11601] = 8'h04 ;
            rom[11602] = 8'heb ;
            rom[11603] = 8'h25 ;
            rom[11604] = 8'hc6 ;
            rom[11605] = 8'h07 ;
            rom[11606] = 8'h12 ;
            rom[11607] = 8'h20 ;
            rom[11608] = 8'h03 ;
            rom[11609] = 8'h0c ;
            rom[11610] = 8'h00 ;
            rom[11611] = 8'h26 ;
            rom[11612] = 8'hed ;
            rom[11613] = 8'hcd ;
            rom[11614] = 8'hf0 ;
            rom[11615] = 8'h0c ;
            rom[11616] = 8'h10 ;
            rom[11617] = 8'h1c ;
            rom[11618] = 8'h04 ;
            rom[11619] = 8'he8 ;
            rom[11620] = 8'he1 ;
            rom[11621] = 8'h08 ;
            rom[11622] = 8'h12 ;
            rom[11623] = 8'he4 ;
            rom[11624] = 8'he5 ;
            rom[11625] = 8'h15 ;
            rom[11626] = 8'hea ;
            rom[11627] = 8'hed ;
            rom[11628] = 8'hfd ;
            rom[11629] = 8'hfa ;
            rom[11630] = 8'h16 ;
            rom[11631] = 8'h09 ;
            rom[11632] = 8'h04 ;
            rom[11633] = 8'he7 ;
            rom[11634] = 8'h19 ;
            rom[11635] = 8'hf2 ;
            rom[11636] = 8'h01 ;
            rom[11637] = 8'hee ;
            rom[11638] = 8'h0e ;
            rom[11639] = 8'h07 ;
            rom[11640] = 8'h13 ;
            rom[11641] = 8'he4 ;
            rom[11642] = 8'h02 ;
            rom[11643] = 8'he5 ;
            rom[11644] = 8'h00 ;
            rom[11645] = 8'h18 ;
            rom[11646] = 8'h0a ;
            rom[11647] = 8'hfe ;
            rom[11648] = 8'h1c ;
            rom[11649] = 8'he8 ;
            rom[11650] = 8'hf5 ;
            rom[11651] = 8'hcf ;
            rom[11652] = 8'he7 ;
            rom[11653] = 8'h0a ;
            rom[11654] = 8'h02 ;
            rom[11655] = 8'hf4 ;
            rom[11656] = 8'h02 ;
            rom[11657] = 8'hfd ;
            rom[11658] = 8'hee ;
            rom[11659] = 8'h06 ;
            rom[11660] = 8'h10 ;
            rom[11661] = 8'he5 ;
            rom[11662] = 8'hdc ;
            rom[11663] = 8'h07 ;
            rom[11664] = 8'he5 ;
            rom[11665] = 8'hf8 ;
            rom[11666] = 8'hf8 ;
            rom[11667] = 8'he2 ;
            rom[11668] = 8'hf7 ;
            rom[11669] = 8'hf7 ;
            rom[11670] = 8'h24 ;
            rom[11671] = 8'h20 ;
            rom[11672] = 8'hd8 ;
            rom[11673] = 8'heb ;
            rom[11674] = 8'hff ;
            rom[11675] = 8'hf2 ;
            rom[11676] = 8'h09 ;
            rom[11677] = 8'hf4 ;
            rom[11678] = 8'hea ;
            rom[11679] = 8'h10 ;
            rom[11680] = 8'h02 ;
            rom[11681] = 8'h15 ;
            rom[11682] = 8'hc0 ;
            rom[11683] = 8'hfc ;
            rom[11684] = 8'hee ;
            rom[11685] = 8'h10 ;
            rom[11686] = 8'h04 ;
            rom[11687] = 8'h1d ;
            rom[11688] = 8'hbe ;
            rom[11689] = 8'hfc ;
            rom[11690] = 8'h14 ;
            rom[11691] = 8'hd5 ;
            rom[11692] = 8'he3 ;
            rom[11693] = 8'h0d ;
            rom[11694] = 8'hf8 ;
            rom[11695] = 8'he9 ;
            rom[11696] = 8'h03 ;
            rom[11697] = 8'hb9 ;
            rom[11698] = 8'hee ;
            rom[11699] = 8'hfc ;
            rom[11700] = 8'he9 ;
            rom[11701] = 8'hf6 ;
            rom[11702] = 8'hd0 ;
            rom[11703] = 8'hf3 ;
            rom[11704] = 8'h00 ;
            rom[11705] = 8'h15 ;
            rom[11706] = 8'h12 ;
            rom[11707] = 8'he6 ;
            rom[11708] = 8'h0a ;
            rom[11709] = 8'h0d ;
            rom[11710] = 8'h00 ;
            rom[11711] = 8'hf1 ;
            rom[11712] = 8'h0e ;
            rom[11713] = 8'hd7 ;
            rom[11714] = 8'h2f ;
            rom[11715] = 8'hee ;
            rom[11716] = 8'he9 ;
            rom[11717] = 8'hf2 ;
            rom[11718] = 8'hec ;
            rom[11719] = 8'h0f ;
            rom[11720] = 8'hf7 ;
            rom[11721] = 8'h01 ;
            rom[11722] = 8'h16 ;
            rom[11723] = 8'h22 ;
            rom[11724] = 8'hd6 ;
            rom[11725] = 8'h03 ;
            rom[11726] = 8'h27 ;
            rom[11727] = 8'h17 ;
            rom[11728] = 8'h02 ;
            rom[11729] = 8'hff ;
            rom[11730] = 8'h07 ;
            rom[11731] = 8'h10 ;
            rom[11732] = 8'hc9 ;
            rom[11733] = 8'h16 ;
            rom[11734] = 8'hd6 ;
            rom[11735] = 8'h10 ;
            rom[11736] = 8'h20 ;
            rom[11737] = 8'h12 ;
            rom[11738] = 8'hec ;
            rom[11739] = 8'h23 ;
            rom[11740] = 8'he3 ;
            rom[11741] = 8'he1 ;
            rom[11742] = 8'hd8 ;
            rom[11743] = 8'heb ;
            rom[11744] = 8'h00 ;
            rom[11745] = 8'h02 ;
            rom[11746] = 8'hda ;
            rom[11747] = 8'hfe ;
            rom[11748] = 8'hf7 ;
            rom[11749] = 8'h02 ;
            rom[11750] = 8'h11 ;
            rom[11751] = 8'h01 ;
            rom[11752] = 8'he6 ;
            rom[11753] = 8'h05 ;
            rom[11754] = 8'h14 ;
            rom[11755] = 8'he1 ;
            rom[11756] = 8'h03 ;
            rom[11757] = 8'hf4 ;
            rom[11758] = 8'h13 ;
            rom[11759] = 8'hfc ;
            rom[11760] = 8'he4 ;
            rom[11761] = 8'hfd ;
            rom[11762] = 8'h18 ;
            rom[11763] = 8'h0f ;
            rom[11764] = 8'h06 ;
            rom[11765] = 8'hfe ;
            rom[11766] = 8'h01 ;
            rom[11767] = 8'hfe ;
            rom[11768] = 8'h1d ;
            rom[11769] = 8'hca ;
            rom[11770] = 8'h10 ;
            rom[11771] = 8'hfb ;
            rom[11772] = 8'h14 ;
            rom[11773] = 8'h20 ;
            rom[11774] = 8'h13 ;
            rom[11775] = 8'h01 ;
            rom[11776] = 8'h0c ;
            rom[11777] = 8'hda ;
            rom[11778] = 8'hd1 ;
            rom[11779] = 8'hdf ;
            rom[11780] = 8'hc9 ;
            rom[11781] = 8'h04 ;
            rom[11782] = 8'h0a ;
            rom[11783] = 8'h0c ;
            rom[11784] = 8'h1b ;
            rom[11785] = 8'h26 ;
            rom[11786] = 8'hf0 ;
            rom[11787] = 8'hd2 ;
            rom[11788] = 8'h06 ;
            rom[11789] = 8'h07 ;
            rom[11790] = 8'hec ;
            rom[11791] = 8'h08 ;
            rom[11792] = 8'hff ;
            rom[11793] = 8'h10 ;
            rom[11794] = 8'h21 ;
            rom[11795] = 8'h05 ;
            rom[11796] = 8'hde ;
            rom[11797] = 8'hfe ;
            rom[11798] = 8'h10 ;
            rom[11799] = 8'h21 ;
            rom[11800] = 8'he3 ;
            rom[11801] = 8'h25 ;
            rom[11802] = 8'hed ;
            rom[11803] = 8'h11 ;
            rom[11804] = 8'hf4 ;
            rom[11805] = 8'hf1 ;
            rom[11806] = 8'hff ;
            rom[11807] = 8'he4 ;
            rom[11808] = 8'hf9 ;
            rom[11809] = 8'hf5 ;
            rom[11810] = 8'hce ;
            rom[11811] = 8'h1b ;
            rom[11812] = 8'h00 ;
            rom[11813] = 8'hea ;
            rom[11814] = 8'heb ;
            rom[11815] = 8'h01 ;
            rom[11816] = 8'h00 ;
            rom[11817] = 8'h00 ;
            rom[11818] = 8'h05 ;
            rom[11819] = 8'hf9 ;
            rom[11820] = 8'h06 ;
            rom[11821] = 8'hda ;
            rom[11822] = 8'h06 ;
            rom[11823] = 8'h0d ;
            rom[11824] = 8'hff ;
            rom[11825] = 8'he7 ;
            rom[11826] = 8'hf5 ;
            rom[11827] = 8'he5 ;
            rom[11828] = 8'h00 ;
            rom[11829] = 8'h05 ;
            rom[11830] = 8'he3 ;
            rom[11831] = 8'hcc ;
            rom[11832] = 8'hf2 ;
            rom[11833] = 8'hec ;
            rom[11834] = 8'hf4 ;
            rom[11835] = 8'h0d ;
            rom[11836] = 8'h14 ;
            rom[11837] = 8'h04 ;
            rom[11838] = 8'he3 ;
            rom[11839] = 8'hf1 ;
            rom[11840] = 8'h03 ;
            rom[11841] = 8'h13 ;
            rom[11842] = 8'hf4 ;
            rom[11843] = 8'heb ;
            rom[11844] = 8'hd6 ;
            rom[11845] = 8'hff ;
            rom[11846] = 8'h0e ;
            rom[11847] = 8'h05 ;
            rom[11848] = 8'he7 ;
            rom[11849] = 8'hf9 ;
            rom[11850] = 8'hc9 ;
            rom[11851] = 8'hef ;
            rom[11852] = 8'he6 ;
            rom[11853] = 8'h07 ;
            rom[11854] = 8'he7 ;
            rom[11855] = 8'h03 ;
            rom[11856] = 8'hd6 ;
            rom[11857] = 8'he5 ;
            rom[11858] = 8'h0c ;
            rom[11859] = 8'heb ;
            rom[11860] = 8'hbf ;
            rom[11861] = 8'hfb ;
            rom[11862] = 8'hfb ;
            rom[11863] = 8'h07 ;
            rom[11864] = 8'hf0 ;
            rom[11865] = 8'h01 ;
            rom[11866] = 8'hfe ;
            rom[11867] = 8'h07 ;
            rom[11868] = 8'hff ;
            rom[11869] = 8'h00 ;
            rom[11870] = 8'h0a ;
            rom[11871] = 8'hc1 ;
            rom[11872] = 8'hf7 ;
            rom[11873] = 8'hdf ;
            rom[11874] = 8'h08 ;
            rom[11875] = 8'hde ;
            rom[11876] = 8'hea ;
            rom[11877] = 8'h11 ;
            rom[11878] = 8'he1 ;
            rom[11879] = 8'hfb ;
            rom[11880] = 8'hfd ;
            rom[11881] = 8'h00 ;
            rom[11882] = 8'hf5 ;
            rom[11883] = 8'hd1 ;
            rom[11884] = 8'hf2 ;
            rom[11885] = 8'hfd ;
            rom[11886] = 8'heb ;
            rom[11887] = 8'h16 ;
            rom[11888] = 8'h04 ;
            rom[11889] = 8'hf8 ;
            rom[11890] = 8'hf2 ;
            rom[11891] = 8'hfd ;
            rom[11892] = 8'hf7 ;
            rom[11893] = 8'hf0 ;
            rom[11894] = 8'he2 ;
            rom[11895] = 8'hf3 ;
            rom[11896] = 8'h07 ;
            rom[11897] = 8'h0d ;
            rom[11898] = 8'hf5 ;
            rom[11899] = 8'he5 ;
            rom[11900] = 8'h06 ;
            rom[11901] = 8'h09 ;
            rom[11902] = 8'h0f ;
            rom[11903] = 8'h07 ;
            rom[11904] = 8'h0c ;
            rom[11905] = 8'hf6 ;
            rom[11906] = 8'h00 ;
            rom[11907] = 8'hc4 ;
            rom[11908] = 8'ha3 ;
            rom[11909] = 8'h05 ;
            rom[11910] = 8'hed ;
            rom[11911] = 8'h17 ;
            rom[11912] = 8'heb ;
            rom[11913] = 8'hed ;
            rom[11914] = 8'hfa ;
            rom[11915] = 8'hf5 ;
            rom[11916] = 8'h06 ;
            rom[11917] = 8'hfb ;
            rom[11918] = 8'hff ;
            rom[11919] = 8'hfb ;
            rom[11920] = 8'hcd ;
            rom[11921] = 8'hfb ;
            rom[11922] = 8'h0c ;
            rom[11923] = 8'hd8 ;
            rom[11924] = 8'h9a ;
            rom[11925] = 8'h03 ;
            rom[11926] = 8'hfd ;
            rom[11927] = 8'h2c ;
            rom[11928] = 8'hf7 ;
            rom[11929] = 8'hdd ;
            rom[11930] = 8'h11 ;
            rom[11931] = 8'h01 ;
            rom[11932] = 8'hfd ;
            rom[11933] = 8'he3 ;
            rom[11934] = 8'h11 ;
            rom[11935] = 8'hf1 ;
            rom[11936] = 8'h17 ;
            rom[11937] = 8'hd7 ;
            rom[11938] = 8'h03 ;
            rom[11939] = 8'hfd ;
            rom[11940] = 8'hf1 ;
            rom[11941] = 8'hf7 ;
            rom[11942] = 8'h05 ;
            rom[11943] = 8'h07 ;
            rom[11944] = 8'heb ;
            rom[11945] = 8'h0a ;
            rom[11946] = 8'heb ;
            rom[11947] = 8'he1 ;
            rom[11948] = 8'hf7 ;
            rom[11949] = 8'h01 ;
            rom[11950] = 8'hfa ;
            rom[11951] = 8'hf6 ;
            rom[11952] = 8'h1b ;
            rom[11953] = 8'hdc ;
            rom[11954] = 8'hed ;
            rom[11955] = 8'h0c ;
            rom[11956] = 8'h0b ;
            rom[11957] = 8'he6 ;
            rom[11958] = 8'hf0 ;
            rom[11959] = 8'hf0 ;
            rom[11960] = 8'h11 ;
            rom[11961] = 8'h0d ;
            rom[11962] = 8'h02 ;
            rom[11963] = 8'he9 ;
            rom[11964] = 8'h0b ;
            rom[11965] = 8'hf4 ;
            rom[11966] = 8'h01 ;
            rom[11967] = 8'h0f ;
            rom[11968] = 8'h0a ;
            rom[11969] = 8'h01 ;
            rom[11970] = 8'h14 ;
            rom[11971] = 8'hee ;
            rom[11972] = 8'hde ;
            rom[11973] = 8'he7 ;
            rom[11974] = 8'he2 ;
            rom[11975] = 8'h11 ;
            rom[11976] = 8'hed ;
            rom[11977] = 8'h10 ;
            rom[11978] = 8'he0 ;
            rom[11979] = 8'h1d ;
            rom[11980] = 8'hed ;
            rom[11981] = 8'hfa ;
            rom[11982] = 8'h0f ;
            rom[11983] = 8'h19 ;
            rom[11984] = 8'hf3 ;
            rom[11985] = 8'hf6 ;
            rom[11986] = 8'h06 ;
            rom[11987] = 8'h12 ;
            rom[11988] = 8'hb0 ;
            rom[11989] = 8'h06 ;
            rom[11990] = 8'hf9 ;
            rom[11991] = 8'h09 ;
            rom[11992] = 8'h01 ;
            rom[11993] = 8'h0c ;
            rom[11994] = 8'hed ;
            rom[11995] = 8'h1e ;
            rom[11996] = 8'hf1 ;
            rom[11997] = 8'hd5 ;
            rom[11998] = 8'hda ;
            rom[11999] = 8'hd3 ;
            rom[12000] = 8'h0f ;
            rom[12001] = 8'hd5 ;
            rom[12002] = 8'hef ;
            rom[12003] = 8'he6 ;
            rom[12004] = 8'hf2 ;
            rom[12005] = 8'he4 ;
            rom[12006] = 8'h08 ;
            rom[12007] = 8'hf6 ;
            rom[12008] = 8'heb ;
            rom[12009] = 8'hfd ;
            rom[12010] = 8'h01 ;
            rom[12011] = 8'hdc ;
            rom[12012] = 8'hfc ;
            rom[12013] = 8'hfe ;
            rom[12014] = 8'hee ;
            rom[12015] = 8'h02 ;
            rom[12016] = 8'h0e ;
            rom[12017] = 8'he5 ;
            rom[12018] = 8'hf1 ;
            rom[12019] = 8'h12 ;
            rom[12020] = 8'h03 ;
            rom[12021] = 8'hfc ;
            rom[12022] = 8'hf9 ;
            rom[12023] = 8'hff ;
            rom[12024] = 8'h0f ;
            rom[12025] = 8'hef ;
            rom[12026] = 8'h10 ;
            rom[12027] = 8'hfc ;
            rom[12028] = 8'h1f ;
            rom[12029] = 8'h16 ;
            rom[12030] = 8'h08 ;
            rom[12031] = 8'hdc ;
            rom[12032] = 8'h15 ;
            rom[12033] = 8'hf3 ;
            rom[12034] = 8'h22 ;
            rom[12035] = 8'h0b ;
            rom[12036] = 8'hda ;
            rom[12037] = 8'he0 ;
            rom[12038] = 8'he3 ;
            rom[12039] = 8'hf7 ;
            rom[12040] = 8'h07 ;
            rom[12041] = 8'he4 ;
            rom[12042] = 8'hfd ;
            rom[12043] = 8'h1a ;
            rom[12044] = 8'h06 ;
            rom[12045] = 8'hf9 ;
            rom[12046] = 8'hf3 ;
            rom[12047] = 8'h19 ;
            rom[12048] = 8'hf8 ;
            rom[12049] = 8'h18 ;
            rom[12050] = 8'h06 ;
            rom[12051] = 8'h0e ;
            rom[12052] = 8'he7 ;
            rom[12053] = 8'h1a ;
            rom[12054] = 8'h10 ;
            rom[12055] = 8'hfc ;
            rom[12056] = 8'h03 ;
            rom[12057] = 8'h09 ;
            rom[12058] = 8'hf5 ;
            rom[12059] = 8'hfa ;
            rom[12060] = 8'hf3 ;
            rom[12061] = 8'hfb ;
            rom[12062] = 8'hc2 ;
            rom[12063] = 8'hf9 ;
            rom[12064] = 8'hff ;
            rom[12065] = 8'h0a ;
            rom[12066] = 8'hfb ;
            rom[12067] = 8'h10 ;
            rom[12068] = 8'hf9 ;
            rom[12069] = 8'hfe ;
            rom[12070] = 8'h1e ;
            rom[12071] = 8'he0 ;
            rom[12072] = 8'he6 ;
            rom[12073] = 8'h01 ;
            rom[12074] = 8'h06 ;
            rom[12075] = 8'hf8 ;
            rom[12076] = 8'h04 ;
            rom[12077] = 8'hd1 ;
            rom[12078] = 8'h17 ;
            rom[12079] = 8'hef ;
            rom[12080] = 8'h16 ;
            rom[12081] = 8'hef ;
            rom[12082] = 8'h1c ;
            rom[12083] = 8'he7 ;
            rom[12084] = 8'h14 ;
            rom[12085] = 8'he7 ;
            rom[12086] = 8'hf6 ;
            rom[12087] = 8'hee ;
            rom[12088] = 8'hd0 ;
            rom[12089] = 8'he6 ;
            rom[12090] = 8'h21 ;
            rom[12091] = 8'hd9 ;
            rom[12092] = 8'h06 ;
            rom[12093] = 8'h1c ;
            rom[12094] = 8'h03 ;
            rom[12095] = 8'he1 ;
            rom[12096] = 8'h01 ;
            rom[12097] = 8'hf5 ;
            rom[12098] = 8'he4 ;
            rom[12099] = 8'hd8 ;
            rom[12100] = 8'h0d ;
            rom[12101] = 8'hfe ;
            rom[12102] = 8'h02 ;
            rom[12103] = 8'hdd ;
            rom[12104] = 8'h1f ;
            rom[12105] = 8'h12 ;
            rom[12106] = 8'h06 ;
            rom[12107] = 8'h08 ;
            rom[12108] = 8'h05 ;
            rom[12109] = 8'h1b ;
            rom[12110] = 8'h08 ;
            rom[12111] = 8'hda ;
            rom[12112] = 8'h18 ;
            rom[12113] = 8'hec ;
            rom[12114] = 8'h02 ;
            rom[12115] = 8'h05 ;
            rom[12116] = 8'hda ;
            rom[12117] = 8'he7 ;
            rom[12118] = 8'hdf ;
            rom[12119] = 8'h00 ;
            rom[12120] = 8'h08 ;
            rom[12121] = 8'he4 ;
            rom[12122] = 8'hf0 ;
            rom[12123] = 8'h03 ;
            rom[12124] = 8'h00 ;
            rom[12125] = 8'h0b ;
            rom[12126] = 8'he6 ;
            rom[12127] = 8'h01 ;
            rom[12128] = 8'h13 ;
            rom[12129] = 8'h07 ;
            rom[12130] = 8'h16 ;
            rom[12131] = 8'hf0 ;
            rom[12132] = 8'h15 ;
            rom[12133] = 8'h11 ;
            rom[12134] = 8'hf1 ;
            rom[12135] = 8'hc2 ;
            rom[12136] = 8'h02 ;
            rom[12137] = 8'hfb ;
            rom[12138] = 8'hfd ;
            rom[12139] = 8'hf9 ;
            rom[12140] = 8'h0d ;
            rom[12141] = 8'hfa ;
            rom[12142] = 8'hfc ;
            rom[12143] = 8'he4 ;
            rom[12144] = 8'hee ;
            rom[12145] = 8'hee ;
            rom[12146] = 8'hdf ;
            rom[12147] = 8'h1b ;
            rom[12148] = 8'hf1 ;
            rom[12149] = 8'hfc ;
            rom[12150] = 8'h1c ;
            rom[12151] = 8'he6 ;
            rom[12152] = 8'h13 ;
            rom[12153] = 8'hf9 ;
            rom[12154] = 8'hde ;
            rom[12155] = 8'h1d ;
            rom[12156] = 8'hfb ;
            rom[12157] = 8'hd7 ;
            rom[12158] = 8'h06 ;
            rom[12159] = 8'h00 ;
            rom[12160] = 8'h0b ;
            rom[12161] = 8'h1b ;
            rom[12162] = 8'hec ;
            rom[12163] = 8'hde ;
            rom[12164] = 8'hd8 ;
            rom[12165] = 8'hfa ;
            rom[12166] = 8'h0a ;
            rom[12167] = 8'hc4 ;
            rom[12168] = 8'h05 ;
            rom[12169] = 8'h1b ;
            rom[12170] = 8'hfb ;
            rom[12171] = 8'hd4 ;
            rom[12172] = 8'he3 ;
            rom[12173] = 8'hf1 ;
            rom[12174] = 8'hf8 ;
            rom[12175] = 8'hee ;
            rom[12176] = 8'h07 ;
            rom[12177] = 8'h11 ;
            rom[12178] = 8'hd7 ;
            rom[12179] = 8'hf2 ;
            rom[12180] = 8'h03 ;
            rom[12181] = 8'hef ;
            rom[12182] = 8'h06 ;
            rom[12183] = 8'hf6 ;
            rom[12184] = 8'hc8 ;
            rom[12185] = 8'hec ;
            rom[12186] = 8'hfa ;
            rom[12187] = 8'h1a ;
            rom[12188] = 8'h1c ;
            rom[12189] = 8'h07 ;
            rom[12190] = 8'hfd ;
            rom[12191] = 8'h1c ;
            rom[12192] = 8'hf3 ;
            rom[12193] = 8'h04 ;
            rom[12194] = 8'hf5 ;
            rom[12195] = 8'h11 ;
            rom[12196] = 8'h08 ;
            rom[12197] = 8'hed ;
            rom[12198] = 8'hb6 ;
            rom[12199] = 8'h0a ;
            rom[12200] = 8'hf9 ;
            rom[12201] = 8'he5 ;
            rom[12202] = 8'hf3 ;
            rom[12203] = 8'h18 ;
            rom[12204] = 8'hfd ;
            rom[12205] = 8'he9 ;
            rom[12206] = 8'heb ;
            rom[12207] = 8'he4 ;
            rom[12208] = 8'hfe ;
            rom[12209] = 8'hec ;
            rom[12210] = 8'h10 ;
            rom[12211] = 8'hd4 ;
            rom[12212] = 8'h00 ;
            rom[12213] = 8'hfc ;
            rom[12214] = 8'he5 ;
            rom[12215] = 8'hf5 ;
            rom[12216] = 8'hfd ;
            rom[12217] = 8'h07 ;
            rom[12218] = 8'he1 ;
            rom[12219] = 8'hcc ;
            rom[12220] = 8'hee ;
            rom[12221] = 8'h08 ;
            rom[12222] = 8'h03 ;
            rom[12223] = 8'hea ;
            rom[12224] = 8'hfc ;
            rom[12225] = 8'hd4 ;
            rom[12226] = 8'h1a ;
            rom[12227] = 8'h18 ;
            rom[12228] = 8'h06 ;
            rom[12229] = 8'h10 ;
            rom[12230] = 8'h00 ;
            rom[12231] = 8'hfd ;
            rom[12232] = 8'h01 ;
            rom[12233] = 8'hef ;
            rom[12234] = 8'h2b ;
            rom[12235] = 8'h2e ;
            rom[12236] = 8'h2a ;
            rom[12237] = 8'h05 ;
            rom[12238] = 8'h18 ;
            rom[12239] = 8'hdd ;
            rom[12240] = 8'hf8 ;
            rom[12241] = 8'h06 ;
            rom[12242] = 8'h02 ;
            rom[12243] = 8'h14 ;
            rom[12244] = 8'hde ;
            rom[12245] = 8'hf3 ;
            rom[12246] = 8'hfd ;
            rom[12247] = 8'hfc ;
            rom[12248] = 8'h10 ;
            rom[12249] = 8'h08 ;
            rom[12250] = 8'he3 ;
            rom[12251] = 8'h12 ;
            rom[12252] = 8'hfe ;
            rom[12253] = 8'hee ;
            rom[12254] = 8'h08 ;
            rom[12255] = 8'h00 ;
            rom[12256] = 8'h01 ;
            rom[12257] = 8'h00 ;
            rom[12258] = 8'h0e ;
            rom[12259] = 8'h03 ;
            rom[12260] = 8'h20 ;
            rom[12261] = 8'h10 ;
            rom[12262] = 8'h0c ;
            rom[12263] = 8'hcc ;
            rom[12264] = 8'hf0 ;
            rom[12265] = 8'hf3 ;
            rom[12266] = 8'hef ;
            rom[12267] = 8'h07 ;
            rom[12268] = 8'h04 ;
            rom[12269] = 8'hfe ;
            rom[12270] = 8'hf7 ;
            rom[12271] = 8'hf2 ;
            rom[12272] = 8'hd0 ;
            rom[12273] = 8'hf7 ;
            rom[12274] = 8'hea ;
            rom[12275] = 8'h15 ;
            rom[12276] = 8'he9 ;
            rom[12277] = 8'hf8 ;
            rom[12278] = 8'h1e ;
            rom[12279] = 8'h13 ;
            rom[12280] = 8'h24 ;
            rom[12281] = 8'hf2 ;
            rom[12282] = 8'h19 ;
            rom[12283] = 8'h02 ;
            rom[12284] = 8'h06 ;
            rom[12285] = 8'he6 ;
            rom[12286] = 8'h22 ;
            rom[12287] = 8'h16 ;
            rom[12288] = 8'h14 ;
            rom[12289] = 8'hd8 ;
            rom[12290] = 8'hf5 ;
            rom[12291] = 8'hf8 ;
            rom[12292] = 8'h25 ;
            rom[12293] = 8'h07 ;
            rom[12294] = 8'hfe ;
            rom[12295] = 8'he7 ;
            rom[12296] = 8'hfc ;
            rom[12297] = 8'h09 ;
            rom[12298] = 8'hfe ;
            rom[12299] = 8'h18 ;
            rom[12300] = 8'hd8 ;
            rom[12301] = 8'hf3 ;
            rom[12302] = 8'he5 ;
            rom[12303] = 8'hf2 ;
            rom[12304] = 8'h0d ;
            rom[12305] = 8'hff ;
            rom[12306] = 8'h07 ;
            rom[12307] = 8'h09 ;
            rom[12308] = 8'h04 ;
            rom[12309] = 8'h05 ;
            rom[12310] = 8'hd1 ;
            rom[12311] = 8'hfe ;
            rom[12312] = 8'hec ;
            rom[12313] = 8'hf5 ;
            rom[12314] = 8'h06 ;
            rom[12315] = 8'hd6 ;
            rom[12316] = 8'h06 ;
            rom[12317] = 8'hed ;
            rom[12318] = 8'hf1 ;
            rom[12319] = 8'hea ;
            rom[12320] = 8'hf7 ;
            rom[12321] = 8'hf0 ;
            rom[12322] = 8'h01 ;
            rom[12323] = 8'h00 ;
            rom[12324] = 8'he6 ;
            rom[12325] = 8'h18 ;
            rom[12326] = 8'hc5 ;
            rom[12327] = 8'hf7 ;
            rom[12328] = 8'h03 ;
            rom[12329] = 8'h01 ;
            rom[12330] = 8'hfb ;
            rom[12331] = 8'hf4 ;
            rom[12332] = 8'h00 ;
            rom[12333] = 8'h02 ;
            rom[12334] = 8'h0c ;
            rom[12335] = 8'hff ;
            rom[12336] = 8'hde ;
            rom[12337] = 8'h1a ;
            rom[12338] = 8'hfd ;
            rom[12339] = 8'he0 ;
            rom[12340] = 8'hf8 ;
            rom[12341] = 8'he9 ;
            rom[12342] = 8'he3 ;
            rom[12343] = 8'h1e ;
            rom[12344] = 8'hde ;
            rom[12345] = 8'hf3 ;
            rom[12346] = 8'h00 ;
            rom[12347] = 8'h06 ;
            rom[12348] = 8'he5 ;
            rom[12349] = 8'h06 ;
            rom[12350] = 8'hde ;
            rom[12351] = 8'hf8 ;
            rom[12352] = 8'h07 ;
            rom[12353] = 8'hfa ;
            rom[12354] = 8'hff ;
            rom[12355] = 8'h0e ;
            rom[12356] = 8'h13 ;
            rom[12357] = 8'h10 ;
            rom[12358] = 8'hde ;
            rom[12359] = 8'he6 ;
            rom[12360] = 8'h05 ;
            rom[12361] = 8'h17 ;
            rom[12362] = 8'h07 ;
            rom[12363] = 8'hfe ;
            rom[12364] = 8'h0f ;
            rom[12365] = 8'h18 ;
            rom[12366] = 8'hf2 ;
            rom[12367] = 8'hde ;
            rom[12368] = 8'hee ;
            rom[12369] = 8'h0e ;
            rom[12370] = 8'hf0 ;
            rom[12371] = 8'h08 ;
            rom[12372] = 8'h09 ;
            rom[12373] = 8'hf7 ;
            rom[12374] = 8'h10 ;
            rom[12375] = 8'h0c ;
            rom[12376] = 8'h02 ;
            rom[12377] = 8'hca ;
            rom[12378] = 8'h09 ;
            rom[12379] = 8'hfb ;
            rom[12380] = 8'h0b ;
            rom[12381] = 8'h1a ;
            rom[12382] = 8'h18 ;
            rom[12383] = 8'h01 ;
            rom[12384] = 8'hd0 ;
            rom[12385] = 8'h0a ;
            rom[12386] = 8'h04 ;
            rom[12387] = 8'h05 ;
            rom[12388] = 8'hf4 ;
            rom[12389] = 8'h00 ;
            rom[12390] = 8'hfd ;
            rom[12391] = 8'hf5 ;
            rom[12392] = 8'h0b ;
            rom[12393] = 8'hfe ;
            rom[12394] = 8'hf5 ;
            rom[12395] = 8'h03 ;
            rom[12396] = 8'h14 ;
            rom[12397] = 8'h0c ;
            rom[12398] = 8'h04 ;
            rom[12399] = 8'h12 ;
            rom[12400] = 8'he6 ;
            rom[12401] = 8'hdd ;
            rom[12402] = 8'h19 ;
            rom[12403] = 8'hc5 ;
            rom[12404] = 8'h15 ;
            rom[12405] = 8'h1e ;
            rom[12406] = 8'hef ;
            rom[12407] = 8'hfd ;
            rom[12408] = 8'h0a ;
            rom[12409] = 8'h03 ;
            rom[12410] = 8'hf6 ;
            rom[12411] = 8'he8 ;
            rom[12412] = 8'hfe ;
            rom[12413] = 8'h10 ;
            rom[12414] = 8'h08 ;
            rom[12415] = 8'hee ;
            rom[12416] = 8'h05 ;
            rom[12417] = 8'h01 ;
            rom[12418] = 8'hf8 ;
            rom[12419] = 8'hf2 ;
            rom[12420] = 8'h02 ;
            rom[12421] = 8'he3 ;
            rom[12422] = 8'hda ;
            rom[12423] = 8'h16 ;
            rom[12424] = 8'h05 ;
            rom[12425] = 8'hd0 ;
            rom[12426] = 8'h00 ;
            rom[12427] = 8'he8 ;
            rom[12428] = 8'h03 ;
            rom[12429] = 8'hf3 ;
            rom[12430] = 8'h06 ;
            rom[12431] = 8'hc9 ;
            rom[12432] = 8'he7 ;
            rom[12433] = 8'hff ;
            rom[12434] = 8'h06 ;
            rom[12435] = 8'h07 ;
            rom[12436] = 8'h0b ;
            rom[12437] = 8'h1e ;
            rom[12438] = 8'h17 ;
            rom[12439] = 8'h10 ;
            rom[12440] = 8'he6 ;
            rom[12441] = 8'h0b ;
            rom[12442] = 8'he4 ;
            rom[12443] = 8'h0c ;
            rom[12444] = 8'hde ;
            rom[12445] = 8'he5 ;
            rom[12446] = 8'hef ;
            rom[12447] = 8'hfe ;
            rom[12448] = 8'hd9 ;
            rom[12449] = 8'hfb ;
            rom[12450] = 8'hfe ;
            rom[12451] = 8'h07 ;
            rom[12452] = 8'h04 ;
            rom[12453] = 8'hf1 ;
            rom[12454] = 8'h04 ;
            rom[12455] = 8'h12 ;
            rom[12456] = 8'he5 ;
            rom[12457] = 8'h0b ;
            rom[12458] = 8'hfe ;
            rom[12459] = 8'hf5 ;
            rom[12460] = 8'he3 ;
            rom[12461] = 8'h05 ;
            rom[12462] = 8'h08 ;
            rom[12463] = 8'hf1 ;
            rom[12464] = 8'hf4 ;
            rom[12465] = 8'h16 ;
            rom[12466] = 8'hf4 ;
            rom[12467] = 8'hdd ;
            rom[12468] = 8'h01 ;
            rom[12469] = 8'h27 ;
            rom[12470] = 8'h0d ;
            rom[12471] = 8'h0c ;
            rom[12472] = 8'hef ;
            rom[12473] = 8'h03 ;
            rom[12474] = 8'h02 ;
            rom[12475] = 8'h0c ;
            rom[12476] = 8'hfd ;
            rom[12477] = 8'hfb ;
            rom[12478] = 8'h0a ;
            rom[12479] = 8'h0e ;
            rom[12480] = 8'hf4 ;
            rom[12481] = 8'h18 ;
            rom[12482] = 8'h02 ;
            rom[12483] = 8'he6 ;
            rom[12484] = 8'h04 ;
            rom[12485] = 8'hec ;
            rom[12486] = 8'hf0 ;
            rom[12487] = 8'h07 ;
            rom[12488] = 8'he3 ;
            rom[12489] = 8'h02 ;
            rom[12490] = 8'hf6 ;
            rom[12491] = 8'h13 ;
            rom[12492] = 8'hf7 ;
            rom[12493] = 8'h19 ;
            rom[12494] = 8'h36 ;
            rom[12495] = 8'hfe ;
            rom[12496] = 8'hf8 ;
            rom[12497] = 8'hd4 ;
            rom[12498] = 8'h16 ;
            rom[12499] = 8'hdb ;
            rom[12500] = 8'hde ;
            rom[12501] = 8'h07 ;
            rom[12502] = 8'hf4 ;
            rom[12503] = 8'he1 ;
            rom[12504] = 8'h19 ;
            rom[12505] = 8'hfc ;
            rom[12506] = 8'h1b ;
            rom[12507] = 8'h0b ;
            rom[12508] = 8'h30 ;
            rom[12509] = 8'he7 ;
            rom[12510] = 8'hfd ;
            rom[12511] = 8'h15 ;
            rom[12512] = 8'h00 ;
            rom[12513] = 8'h29 ;
            rom[12514] = 8'h10 ;
            rom[12515] = 8'h03 ;
            rom[12516] = 8'h21 ;
            rom[12517] = 8'he8 ;
            rom[12518] = 8'hdb ;
            rom[12519] = 8'h0f ;
            rom[12520] = 8'hf7 ;
            rom[12521] = 8'h10 ;
            rom[12522] = 8'h3a ;
            rom[12523] = 8'hf2 ;
            rom[12524] = 8'h00 ;
            rom[12525] = 8'h0a ;
            rom[12526] = 8'h01 ;
            rom[12527] = 8'hcf ;
            rom[12528] = 8'h19 ;
            rom[12529] = 8'h17 ;
            rom[12530] = 8'hfe ;
            rom[12531] = 8'hf1 ;
            rom[12532] = 8'he8 ;
            rom[12533] = 8'heb ;
            rom[12534] = 8'h07 ;
            rom[12535] = 8'h3a ;
            rom[12536] = 8'hf6 ;
            rom[12537] = 8'h05 ;
            rom[12538] = 8'h0d ;
            rom[12539] = 8'hf6 ;
            rom[12540] = 8'hf9 ;
            rom[12541] = 8'h14 ;
            rom[12542] = 8'hf0 ;
            rom[12543] = 8'h08 ;
            rom[12544] = 8'h11 ;
            rom[12545] = 8'hf3 ;
            rom[12546] = 8'h18 ;
            rom[12547] = 8'h31 ;
            rom[12548] = 8'hfd ;
            rom[12549] = 8'hfd ;
            rom[12550] = 8'h09 ;
            rom[12551] = 8'hef ;
            rom[12552] = 8'hfb ;
            rom[12553] = 8'h01 ;
            rom[12554] = 8'h20 ;
            rom[12555] = 8'h17 ;
            rom[12556] = 8'hf4 ;
            rom[12557] = 8'h20 ;
            rom[12558] = 8'hf2 ;
            rom[12559] = 8'h01 ;
            rom[12560] = 8'hc4 ;
            rom[12561] = 8'hbe ;
            rom[12562] = 8'h03 ;
            rom[12563] = 8'h1c ;
            rom[12564] = 8'hf3 ;
            rom[12565] = 8'hea ;
            rom[12566] = 8'hda ;
            rom[12567] = 8'h11 ;
            rom[12568] = 8'h0f ;
            rom[12569] = 8'hf1 ;
            rom[12570] = 8'hd4 ;
            rom[12571] = 8'h03 ;
            rom[12572] = 8'hf9 ;
            rom[12573] = 8'hf2 ;
            rom[12574] = 8'h03 ;
            rom[12575] = 8'he5 ;
            rom[12576] = 8'hf5 ;
            rom[12577] = 8'h0a ;
            rom[12578] = 8'hf0 ;
            rom[12579] = 8'he0 ;
            rom[12580] = 8'h23 ;
            rom[12581] = 8'hfa ;
            rom[12582] = 8'hfc ;
            rom[12583] = 8'hf1 ;
            rom[12584] = 8'h16 ;
            rom[12585] = 8'hd5 ;
            rom[12586] = 8'hef ;
            rom[12587] = 8'h07 ;
            rom[12588] = 8'hd6 ;
            rom[12589] = 8'h05 ;
            rom[12590] = 8'hf8 ;
            rom[12591] = 8'hfc ;
            rom[12592] = 8'he4 ;
            rom[12593] = 8'hff ;
            rom[12594] = 8'h0d ;
            rom[12595] = 8'h00 ;
            rom[12596] = 8'hf9 ;
            rom[12597] = 8'h10 ;
            rom[12598] = 8'hf7 ;
            rom[12599] = 8'hf4 ;
            rom[12600] = 8'hff ;
            rom[12601] = 8'hf1 ;
            rom[12602] = 8'hfa ;
            rom[12603] = 8'h00 ;
            rom[12604] = 8'hf9 ;
            rom[12605] = 8'h03 ;
            rom[12606] = 8'he1 ;
            rom[12607] = 8'hf6 ;
            rom[12608] = 8'h0a ;
            rom[12609] = 8'h13 ;
            rom[12610] = 8'h04 ;
            rom[12611] = 8'h09 ;
            rom[12612] = 8'hf5 ;
            rom[12613] = 8'hfc ;
            rom[12614] = 8'h17 ;
            rom[12615] = 8'h28 ;
            rom[12616] = 8'hfc ;
            rom[12617] = 8'h05 ;
            rom[12618] = 8'h08 ;
            rom[12619] = 8'hdf ;
            rom[12620] = 8'h0a ;
            rom[12621] = 8'h1f ;
            rom[12622] = 8'h18 ;
            rom[12623] = 8'hba ;
            rom[12624] = 8'hd7 ;
            rom[12625] = 8'hf4 ;
            rom[12626] = 8'hf5 ;
            rom[12627] = 8'h03 ;
            rom[12628] = 8'hfa ;
            rom[12629] = 8'hdb ;
            rom[12630] = 8'hd2 ;
            rom[12631] = 8'h13 ;
            rom[12632] = 8'h09 ;
            rom[12633] = 8'hf2 ;
            rom[12634] = 8'hee ;
            rom[12635] = 8'h15 ;
            rom[12636] = 8'h04 ;
            rom[12637] = 8'hf8 ;
            rom[12638] = 8'h07 ;
            rom[12639] = 8'hfd ;
            rom[12640] = 8'hf9 ;
            rom[12641] = 8'h00 ;
            rom[12642] = 8'heb ;
            rom[12643] = 8'h0e ;
            rom[12644] = 8'h1c ;
            rom[12645] = 8'h0c ;
            rom[12646] = 8'hf7 ;
            rom[12647] = 8'h20 ;
            rom[12648] = 8'hfc ;
            rom[12649] = 8'h0b ;
            rom[12650] = 8'hf1 ;
            rom[12651] = 8'h33 ;
            rom[12652] = 8'hf4 ;
            rom[12653] = 8'h0c ;
            rom[12654] = 8'hef ;
            rom[12655] = 8'he2 ;
            rom[12656] = 8'hd7 ;
            rom[12657] = 8'h17 ;
            rom[12658] = 8'h16 ;
            rom[12659] = 8'hf8 ;
            rom[12660] = 8'hd7 ;
            rom[12661] = 8'h08 ;
            rom[12662] = 8'h0f ;
            rom[12663] = 8'h14 ;
            rom[12664] = 8'h08 ;
            rom[12665] = 8'hf5 ;
            rom[12666] = 8'h07 ;
            rom[12667] = 8'h12 ;
            rom[12668] = 8'h0d ;
            rom[12669] = 8'hd2 ;
            rom[12670] = 8'h14 ;
            rom[12671] = 8'hfa ;
            rom[12672] = 8'h0f ;
            rom[12673] = 8'he6 ;
            rom[12674] = 8'hfb ;
            rom[12675] = 8'h07 ;
            rom[12676] = 8'h0b ;
            rom[12677] = 8'hc7 ;
            rom[12678] = 8'hf5 ;
            rom[12679] = 8'hf5 ;
            rom[12680] = 8'he8 ;
            rom[12681] = 8'hda ;
            rom[12682] = 8'hf1 ;
            rom[12683] = 8'h12 ;
            rom[12684] = 8'he9 ;
            rom[12685] = 8'h18 ;
            rom[12686] = 8'h1a ;
            rom[12687] = 8'h08 ;
            rom[12688] = 8'hf0 ;
            rom[12689] = 8'h32 ;
            rom[12690] = 8'h16 ;
            rom[12691] = 8'h12 ;
            rom[12692] = 8'h04 ;
            rom[12693] = 8'h06 ;
            rom[12694] = 8'h15 ;
            rom[12695] = 8'he5 ;
            rom[12696] = 8'hee ;
            rom[12697] = 8'hf5 ;
            rom[12698] = 8'h1b ;
            rom[12699] = 8'h07 ;
            rom[12700] = 8'hd5 ;
            rom[12701] = 8'heb ;
            rom[12702] = 8'h21 ;
            rom[12703] = 8'h1b ;
            rom[12704] = 8'hc2 ;
            rom[12705] = 8'hf5 ;
            rom[12706] = 8'he2 ;
            rom[12707] = 8'h0a ;
            rom[12708] = 8'h03 ;
            rom[12709] = 8'h1d ;
            rom[12710] = 8'hf1 ;
            rom[12711] = 8'h19 ;
            rom[12712] = 8'h02 ;
            rom[12713] = 8'hfa ;
            rom[12714] = 8'h09 ;
            rom[12715] = 8'h02 ;
            rom[12716] = 8'h0e ;
            rom[12717] = 8'hec ;
            rom[12718] = 8'hd3 ;
            rom[12719] = 8'hf9 ;
            rom[12720] = 8'h20 ;
            rom[12721] = 8'h0c ;
            rom[12722] = 8'hbc ;
            rom[12723] = 8'hec ;
            rom[12724] = 8'h02 ;
            rom[12725] = 8'h10 ;
            rom[12726] = 8'h24 ;
            rom[12727] = 8'hff ;
            rom[12728] = 8'hec ;
            rom[12729] = 8'h37 ;
            rom[12730] = 8'heb ;
            rom[12731] = 8'h10 ;
            rom[12732] = 8'he0 ;
            rom[12733] = 8'hf1 ;
            rom[12734] = 8'hfd ;
            rom[12735] = 8'hfd ;
            rom[12736] = 8'h36 ;
            rom[12737] = 8'h0d ;
            rom[12738] = 8'he4 ;
            rom[12739] = 8'hfb ;
            rom[12740] = 8'hf1 ;
            rom[12741] = 8'hf2 ;
            rom[12742] = 8'hc8 ;
            rom[12743] = 8'h1e ;
            rom[12744] = 8'hd6 ;
            rom[12745] = 8'hf8 ;
            rom[12746] = 8'h11 ;
            rom[12747] = 8'hf1 ;
            rom[12748] = 8'hde ;
            rom[12749] = 8'hdd ;
            rom[12750] = 8'h0e ;
            rom[12751] = 8'h00 ;
            rom[12752] = 8'hef ;
            rom[12753] = 8'hfb ;
            rom[12754] = 8'h14 ;
            rom[12755] = 8'h01 ;
            rom[12756] = 8'hf0 ;
            rom[12757] = 8'hfb ;
            rom[12758] = 8'hf1 ;
            rom[12759] = 8'h11 ;
            rom[12760] = 8'h05 ;
            rom[12761] = 8'hfe ;
            rom[12762] = 8'h01 ;
            rom[12763] = 8'hf3 ;
            rom[12764] = 8'hfd ;
            rom[12765] = 8'heb ;
            rom[12766] = 8'h0f ;
            rom[12767] = 8'h03 ;
            rom[12768] = 8'he9 ;
            rom[12769] = 8'hee ;
            rom[12770] = 8'hf5 ;
            rom[12771] = 8'h10 ;
            rom[12772] = 8'hf5 ;
            rom[12773] = 8'h32 ;
            rom[12774] = 8'h20 ;
            rom[12775] = 8'h07 ;
            rom[12776] = 8'hfa ;
            rom[12777] = 8'hf8 ;
            rom[12778] = 8'hf1 ;
            rom[12779] = 8'h12 ;
            rom[12780] = 8'hf1 ;
            rom[12781] = 8'hf0 ;
            rom[12782] = 8'h1b ;
            rom[12783] = 8'hd2 ;
            rom[12784] = 8'h19 ;
            rom[12785] = 8'h04 ;
            rom[12786] = 8'h07 ;
            rom[12787] = 8'he6 ;
            rom[12788] = 8'h09 ;
            rom[12789] = 8'hfe ;
            rom[12790] = 8'hfe ;
            rom[12791] = 8'h0f ;
            rom[12792] = 8'h13 ;
            rom[12793] = 8'hfc ;
            rom[12794] = 8'h18 ;
            rom[12795] = 8'hef ;
            rom[12796] = 8'h0a ;
            rom[12797] = 8'hcd ;
            rom[12798] = 8'hf4 ;
            rom[12799] = 8'hfb ;
            rom[12800] = 8'h0e ;
            rom[12801] = 8'h1b ;
            rom[12802] = 8'h02 ;
            rom[12803] = 8'h0e ;
            rom[12804] = 8'h02 ;
            rom[12805] = 8'h05 ;
            rom[12806] = 8'h1d ;
            rom[12807] = 8'hf4 ;
            rom[12808] = 8'hf4 ;
            rom[12809] = 8'he4 ;
            rom[12810] = 8'h1d ;
            rom[12811] = 8'h13 ;
            rom[12812] = 8'h07 ;
            rom[12813] = 8'h0c ;
            rom[12814] = 8'hf7 ;
            rom[12815] = 8'hf1 ;
            rom[12816] = 8'hdc ;
            rom[12817] = 8'h19 ;
            rom[12818] = 8'hff ;
            rom[12819] = 8'hed ;
            rom[12820] = 8'h02 ;
            rom[12821] = 8'he9 ;
            rom[12822] = 8'h0b ;
            rom[12823] = 8'h00 ;
            rom[12824] = 8'h13 ;
            rom[12825] = 8'hb8 ;
            rom[12826] = 8'h13 ;
            rom[12827] = 8'hf2 ;
            rom[12828] = 8'h13 ;
            rom[12829] = 8'h1c ;
            rom[12830] = 8'h04 ;
            rom[12831] = 8'hf4 ;
            rom[12832] = 8'h0b ;
            rom[12833] = 8'h02 ;
            rom[12834] = 8'h07 ;
            rom[12835] = 8'hd3 ;
            rom[12836] = 8'h19 ;
            rom[12837] = 8'h12 ;
            rom[12838] = 8'h0b ;
            rom[12839] = 8'hfd ;
            rom[12840] = 8'h0f ;
            rom[12841] = 8'hb9 ;
            rom[12842] = 8'hf9 ;
            rom[12843] = 8'h27 ;
            rom[12844] = 8'h14 ;
            rom[12845] = 8'hf5 ;
            rom[12846] = 8'hff ;
            rom[12847] = 8'hfb ;
            rom[12848] = 8'h02 ;
            rom[12849] = 8'hd0 ;
            rom[12850] = 8'h14 ;
            rom[12851] = 8'hea ;
            rom[12852] = 8'h08 ;
            rom[12853] = 8'hfe ;
            rom[12854] = 8'h0b ;
            rom[12855] = 8'h14 ;
            rom[12856] = 8'h16 ;
            rom[12857] = 8'h0f ;
            rom[12858] = 8'h0e ;
            rom[12859] = 8'hf6 ;
            rom[12860] = 8'h07 ;
            rom[12861] = 8'h09 ;
            rom[12862] = 8'h02 ;
            rom[12863] = 8'hfa ;
            rom[12864] = 8'h05 ;
            rom[12865] = 8'h08 ;
            rom[12866] = 8'h00 ;
            rom[12867] = 8'h01 ;
            rom[12868] = 8'hf6 ;
            rom[12869] = 8'h06 ;
            rom[12870] = 8'h0a ;
            rom[12871] = 8'hfd ;
            rom[12872] = 8'hf9 ;
            rom[12873] = 8'hfb ;
            rom[12874] = 8'h11 ;
            rom[12875] = 8'hf7 ;
            rom[12876] = 8'h0e ;
            rom[12877] = 8'h1a ;
            rom[12878] = 8'hf4 ;
            rom[12879] = 8'hca ;
            rom[12880] = 8'he8 ;
            rom[12881] = 8'h02 ;
            rom[12882] = 8'he2 ;
            rom[12883] = 8'hfd ;
            rom[12884] = 8'h0f ;
            rom[12885] = 8'hd7 ;
            rom[12886] = 8'hf7 ;
            rom[12887] = 8'h0a ;
            rom[12888] = 8'h05 ;
            rom[12889] = 8'hce ;
            rom[12890] = 8'he6 ;
            rom[12891] = 8'h0a ;
            rom[12892] = 8'h09 ;
            rom[12893] = 8'h0a ;
            rom[12894] = 8'hfc ;
            rom[12895] = 8'hf7 ;
            rom[12896] = 8'hf8 ;
            rom[12897] = 8'hf9 ;
            rom[12898] = 8'h08 ;
            rom[12899] = 8'hd7 ;
            rom[12900] = 8'hf5 ;
            rom[12901] = 8'h0b ;
            rom[12902] = 8'h05 ;
            rom[12903] = 8'he4 ;
            rom[12904] = 8'h22 ;
            rom[12905] = 8'h02 ;
            rom[12906] = 8'hfa ;
            rom[12907] = 8'h15 ;
            rom[12908] = 8'h1b ;
            rom[12909] = 8'hf4 ;
            rom[12910] = 8'hea ;
            rom[12911] = 8'h13 ;
            rom[12912] = 8'hee ;
            rom[12913] = 8'hfa ;
            rom[12914] = 8'h06 ;
            rom[12915] = 8'hd0 ;
            rom[12916] = 8'hfd ;
            rom[12917] = 8'h06 ;
            rom[12918] = 8'h1e ;
            rom[12919] = 8'h0f ;
            rom[12920] = 8'h11 ;
            rom[12921] = 8'h11 ;
            rom[12922] = 8'hf8 ;
            rom[12923] = 8'he7 ;
            rom[12924] = 8'hf5 ;
            rom[12925] = 8'h11 ;
            rom[12926] = 8'h12 ;
            rom[12927] = 8'hde ;
            rom[12928] = 8'hff ;
            rom[12929] = 8'h13 ;
            rom[12930] = 8'h12 ;
            rom[12931] = 8'h11 ;
            rom[12932] = 8'h08 ;
            rom[12933] = 8'h09 ;
            rom[12934] = 8'h13 ;
            rom[12935] = 8'h08 ;
            rom[12936] = 8'hec ;
            rom[12937] = 8'h14 ;
            rom[12938] = 8'hed ;
            rom[12939] = 8'h08 ;
            rom[12940] = 8'h12 ;
            rom[12941] = 8'hfe ;
            rom[12942] = 8'h19 ;
            rom[12943] = 8'hf7 ;
            rom[12944] = 8'hef ;
            rom[12945] = 8'hfd ;
            rom[12946] = 8'h0e ;
            rom[12947] = 8'h1a ;
            rom[12948] = 8'h02 ;
            rom[12949] = 8'hf7 ;
            rom[12950] = 8'hec ;
            rom[12951] = 8'hfa ;
            rom[12952] = 8'hfc ;
            rom[12953] = 8'h04 ;
            rom[12954] = 8'hea ;
            rom[12955] = 8'he0 ;
            rom[12956] = 8'h01 ;
            rom[12957] = 8'hfe ;
            rom[12958] = 8'h1f ;
            rom[12959] = 8'h15 ;
            rom[12960] = 8'hde ;
            rom[12961] = 8'h00 ;
            rom[12962] = 8'h0a ;
            rom[12963] = 8'he2 ;
            rom[12964] = 8'h0b ;
            rom[12965] = 8'h00 ;
            rom[12966] = 8'h13 ;
            rom[12967] = 8'he7 ;
            rom[12968] = 8'h06 ;
            rom[12969] = 8'h02 ;
            rom[12970] = 8'hd6 ;
            rom[12971] = 8'h17 ;
            rom[12972] = 8'h1a ;
            rom[12973] = 8'h06 ;
            rom[12974] = 8'hec ;
            rom[12975] = 8'h1c ;
            rom[12976] = 8'hf1 ;
            rom[12977] = 8'h21 ;
            rom[12978] = 8'h12 ;
            rom[12979] = 8'hf8 ;
            rom[12980] = 8'he9 ;
            rom[12981] = 8'h05 ;
            rom[12982] = 8'h22 ;
            rom[12983] = 8'h13 ;
            rom[12984] = 8'he2 ;
            rom[12985] = 8'hf4 ;
            rom[12986] = 8'h19 ;
            rom[12987] = 8'h2f ;
            rom[12988] = 8'h03 ;
            rom[12989] = 8'hdf ;
            rom[12990] = 8'h0b ;
            rom[12991] = 8'h19 ;
            rom[12992] = 8'h10 ;
            rom[12993] = 8'hfd ;
            rom[12994] = 8'hfa ;
            rom[12995] = 8'h0f ;
            rom[12996] = 8'h05 ;
            rom[12997] = 8'hfa ;
            rom[12998] = 8'h19 ;
            rom[12999] = 8'h02 ;
            rom[13000] = 8'h08 ;
            rom[13001] = 8'hf9 ;
            rom[13002] = 8'h0c ;
            rom[13003] = 8'hf0 ;
            rom[13004] = 8'h09 ;
            rom[13005] = 8'h0a ;
            rom[13006] = 8'h0c ;
            rom[13007] = 8'hfd ;
            rom[13008] = 8'hf2 ;
            rom[13009] = 8'hfd ;
            rom[13010] = 8'hfd ;
            rom[13011] = 8'hfe ;
            rom[13012] = 8'hf8 ;
            rom[13013] = 8'hf9 ;
            rom[13014] = 8'h02 ;
            rom[13015] = 8'h00 ;
            rom[13016] = 8'hf1 ;
            rom[13017] = 8'h07 ;
            rom[13018] = 8'hd9 ;
            rom[13019] = 8'h20 ;
            rom[13020] = 8'h02 ;
            rom[13021] = 8'h0b ;
            rom[13022] = 8'hfb ;
            rom[13023] = 8'h06 ;
            rom[13024] = 8'h15 ;
            rom[13025] = 8'h03 ;
            rom[13026] = 8'h18 ;
            rom[13027] = 8'h01 ;
            rom[13028] = 8'h04 ;
            rom[13029] = 8'h18 ;
            rom[13030] = 8'hf5 ;
            rom[13031] = 8'hdf ;
            rom[13032] = 8'hf8 ;
            rom[13033] = 8'hee ;
            rom[13034] = 8'h02 ;
            rom[13035] = 8'h05 ;
            rom[13036] = 8'h05 ;
            rom[13037] = 8'h07 ;
            rom[13038] = 8'hf8 ;
            rom[13039] = 8'h1e ;
            rom[13040] = 8'hdd ;
            rom[13041] = 8'h0b ;
            rom[13042] = 8'hfb ;
            rom[13043] = 8'hed ;
            rom[13044] = 8'h15 ;
            rom[13045] = 8'h08 ;
            rom[13046] = 8'h11 ;
            rom[13047] = 8'h05 ;
            rom[13048] = 8'hf7 ;
            rom[13049] = 8'h02 ;
            rom[13050] = 8'h16 ;
            rom[13051] = 8'h02 ;
            rom[13052] = 8'h03 ;
            rom[13053] = 8'h0d ;
            rom[13054] = 8'hf2 ;
            rom[13055] = 8'h01 ;
            rom[13056] = 8'hfe ;
            rom[13057] = 8'hf2 ;
            rom[13058] = 8'h0f ;
            rom[13059] = 8'hf1 ;
            rom[13060] = 8'h0a ;
            rom[13061] = 8'hff ;
            rom[13062] = 8'he8 ;
            rom[13063] = 8'he6 ;
            rom[13064] = 8'he1 ;
            rom[13065] = 8'h0c ;
            rom[13066] = 8'hf3 ;
            rom[13067] = 8'he7 ;
            rom[13068] = 8'h1a ;
            rom[13069] = 8'h0f ;
            rom[13070] = 8'hd8 ;
            rom[13071] = 8'hfa ;
            rom[13072] = 8'hf2 ;
            rom[13073] = 8'h15 ;
            rom[13074] = 8'h08 ;
            rom[13075] = 8'h0a ;
            rom[13076] = 8'h02 ;
            rom[13077] = 8'h0a ;
            rom[13078] = 8'h17 ;
            rom[13079] = 8'h0b ;
            rom[13080] = 8'hfe ;
            rom[13081] = 8'hf3 ;
            rom[13082] = 8'h21 ;
            rom[13083] = 8'hfc ;
            rom[13084] = 8'hcf ;
            rom[13085] = 8'hf3 ;
            rom[13086] = 8'h11 ;
            rom[13087] = 8'h0e ;
            rom[13088] = 8'hdc ;
            rom[13089] = 8'hf4 ;
            rom[13090] = 8'heb ;
            rom[13091] = 8'h0c ;
            rom[13092] = 8'he1 ;
            rom[13093] = 8'h02 ;
            rom[13094] = 8'hec ;
            rom[13095] = 8'h14 ;
            rom[13096] = 8'h10 ;
            rom[13097] = 8'hf5 ;
            rom[13098] = 8'hf8 ;
            rom[13099] = 8'hfe ;
            rom[13100] = 8'h00 ;
            rom[13101] = 8'hec ;
            rom[13102] = 8'he0 ;
            rom[13103] = 8'hdf ;
            rom[13104] = 8'h29 ;
            rom[13105] = 8'h08 ;
            rom[13106] = 8'h0b ;
            rom[13107] = 8'he4 ;
            rom[13108] = 8'h10 ;
            rom[13109] = 8'h07 ;
            rom[13110] = 8'h1a ;
            rom[13111] = 8'h11 ;
            rom[13112] = 8'h20 ;
            rom[13113] = 8'h11 ;
            rom[13114] = 8'hda ;
            rom[13115] = 8'h00 ;
            rom[13116] = 8'hd2 ;
            rom[13117] = 8'h07 ;
            rom[13118] = 8'h0e ;
            rom[13119] = 8'h0e ;
            rom[13120] = 8'h1a ;
            rom[13121] = 8'h0a ;
            rom[13122] = 8'h2e ;
            rom[13123] = 8'h03 ;
            rom[13124] = 8'hee ;
            rom[13125] = 8'h0d ;
            rom[13126] = 8'h1e ;
            rom[13127] = 8'hda ;
            rom[13128] = 8'hd4 ;
            rom[13129] = 8'hf2 ;
            rom[13130] = 8'h13 ;
            rom[13131] = 8'h05 ;
            rom[13132] = 8'hd9 ;
            rom[13133] = 8'h15 ;
            rom[13134] = 8'hea ;
            rom[13135] = 8'he4 ;
            rom[13136] = 8'hef ;
            rom[13137] = 8'hf2 ;
            rom[13138] = 8'h07 ;
            rom[13139] = 8'hd0 ;
            rom[13140] = 8'hcc ;
            rom[13141] = 8'hff ;
            rom[13142] = 8'heb ;
            rom[13143] = 8'hf9 ;
            rom[13144] = 8'hf5 ;
            rom[13145] = 8'h00 ;
            rom[13146] = 8'he3 ;
            rom[13147] = 8'hf1 ;
            rom[13148] = 8'he6 ;
            rom[13149] = 8'h07 ;
            rom[13150] = 8'h1e ;
            rom[13151] = 8'hfc ;
            rom[13152] = 8'h04 ;
            rom[13153] = 8'h03 ;
            rom[13154] = 8'h14 ;
            rom[13155] = 8'h0f ;
            rom[13156] = 8'heb ;
            rom[13157] = 8'hff ;
            rom[13158] = 8'he8 ;
            rom[13159] = 8'h12 ;
            rom[13160] = 8'h0f ;
            rom[13161] = 8'h00 ;
            rom[13162] = 8'h20 ;
            rom[13163] = 8'hf2 ;
            rom[13164] = 8'h0b ;
            rom[13165] = 8'h02 ;
            rom[13166] = 8'h05 ;
            rom[13167] = 8'hb5 ;
            rom[13168] = 8'hff ;
            rom[13169] = 8'h07 ;
            rom[13170] = 8'hff ;
            rom[13171] = 8'h08 ;
            rom[13172] = 8'hbd ;
            rom[13173] = 8'hef ;
            rom[13174] = 8'hdf ;
            rom[13175] = 8'h3e ;
            rom[13176] = 8'he8 ;
            rom[13177] = 8'hfc ;
            rom[13178] = 8'hfa ;
            rom[13179] = 8'h14 ;
            rom[13180] = 8'hed ;
            rom[13181] = 8'h01 ;
            rom[13182] = 8'hef ;
            rom[13183] = 8'h28 ;
            rom[13184] = 8'h0a ;
            rom[13185] = 8'hf0 ;
            rom[13186] = 8'heb ;
            rom[13187] = 8'h06 ;
            rom[13188] = 8'h24 ;
            rom[13189] = 8'hf1 ;
            rom[13190] = 8'hfc ;
            rom[13191] = 8'h0e ;
            rom[13192] = 8'hf7 ;
            rom[13193] = 8'hb1 ;
            rom[13194] = 8'hfe ;
            rom[13195] = 8'hf0 ;
            rom[13196] = 8'h13 ;
            rom[13197] = 8'h2c ;
            rom[13198] = 8'h10 ;
            rom[13199] = 8'hee ;
            rom[13200] = 8'hf9 ;
            rom[13201] = 8'h01 ;
            rom[13202] = 8'hff ;
            rom[13203] = 8'h12 ;
            rom[13204] = 8'h03 ;
            rom[13205] = 8'h02 ;
            rom[13206] = 8'hf5 ;
            rom[13207] = 8'hc0 ;
            rom[13208] = 8'hf1 ;
            rom[13209] = 8'h0e ;
            rom[13210] = 8'h1e ;
            rom[13211] = 8'hea ;
            rom[13212] = 8'he2 ;
            rom[13213] = 8'hf9 ;
            rom[13214] = 8'hea ;
            rom[13215] = 8'h0e ;
            rom[13216] = 8'hf9 ;
            rom[13217] = 8'h08 ;
            rom[13218] = 8'h15 ;
            rom[13219] = 8'hf8 ;
            rom[13220] = 8'h11 ;
            rom[13221] = 8'h0d ;
            rom[13222] = 8'he5 ;
            rom[13223] = 8'h0c ;
            rom[13224] = 8'hf7 ;
            rom[13225] = 8'hfd ;
            rom[13226] = 8'hf9 ;
            rom[13227] = 8'hf4 ;
            rom[13228] = 8'h23 ;
            rom[13229] = 8'h0b ;
            rom[13230] = 8'hff ;
            rom[13231] = 8'hfd ;
            rom[13232] = 8'h0f ;
            rom[13233] = 8'h08 ;
            rom[13234] = 8'h1c ;
            rom[13235] = 8'hfd ;
            rom[13236] = 8'he7 ;
            rom[13237] = 8'h2d ;
            rom[13238] = 8'hfc ;
            rom[13239] = 8'hec ;
            rom[13240] = 8'hfe ;
            rom[13241] = 8'h24 ;
            rom[13242] = 8'h0a ;
            rom[13243] = 8'h04 ;
            rom[13244] = 8'h00 ;
            rom[13245] = 8'hc7 ;
            rom[13246] = 8'hf1 ;
            rom[13247] = 8'he3 ;
            rom[13248] = 8'h01 ;
            rom[13249] = 8'hf7 ;
            rom[13250] = 8'hff ;
            rom[13251] = 8'hf9 ;
            rom[13252] = 8'h06 ;
            rom[13253] = 8'hfd ;
            rom[13254] = 8'hf6 ;
            rom[13255] = 8'h0a ;
            rom[13256] = 8'he1 ;
            rom[13257] = 8'hf9 ;
            rom[13258] = 8'h0c ;
            rom[13259] = 8'hf6 ;
            rom[13260] = 8'h1c ;
            rom[13261] = 8'h19 ;
            rom[13262] = 8'h00 ;
            rom[13263] = 8'hf1 ;
            rom[13264] = 8'hf4 ;
            rom[13265] = 8'he2 ;
            rom[13266] = 8'hf2 ;
            rom[13267] = 8'hee ;
            rom[13268] = 8'h0b ;
            rom[13269] = 8'h13 ;
            rom[13270] = 8'h18 ;
            rom[13271] = 8'hf7 ;
            rom[13272] = 8'he5 ;
            rom[13273] = 8'h18 ;
            rom[13274] = 8'hf5 ;
            rom[13275] = 8'h0d ;
            rom[13276] = 8'hf5 ;
            rom[13277] = 8'h02 ;
            rom[13278] = 8'hf0 ;
            rom[13279] = 8'h04 ;
            rom[13280] = 8'h01 ;
            rom[13281] = 8'hf8 ;
            rom[13282] = 8'h0e ;
            rom[13283] = 8'hf7 ;
            rom[13284] = 8'hd0 ;
            rom[13285] = 8'h0f ;
            rom[13286] = 8'hf4 ;
            rom[13287] = 8'hfd ;
            rom[13288] = 8'h1a ;
            rom[13289] = 8'h11 ;
            rom[13290] = 8'hfa ;
            rom[13291] = 8'hf3 ;
            rom[13292] = 8'hf9 ;
            rom[13293] = 8'h17 ;
            rom[13294] = 8'h05 ;
            rom[13295] = 8'hfc ;
            rom[13296] = 8'hda ;
            rom[13297] = 8'h0e ;
            rom[13298] = 8'hf3 ;
            rom[13299] = 8'hf0 ;
            rom[13300] = 8'h02 ;
            rom[13301] = 8'h25 ;
            rom[13302] = 8'hfc ;
            rom[13303] = 8'h12 ;
            rom[13304] = 8'hf7 ;
            rom[13305] = 8'hf9 ;
            rom[13306] = 8'h0d ;
            rom[13307] = 8'h02 ;
            rom[13308] = 8'hd4 ;
            rom[13309] = 8'h16 ;
            rom[13310] = 8'h1a ;
            rom[13311] = 8'h11 ;
            rom[13312] = 8'he7 ;
            rom[13313] = 8'h06 ;
            rom[13314] = 8'h03 ;
            rom[13315] = 8'h16 ;
            rom[13316] = 8'h1e ;
            rom[13317] = 8'hfc ;
            rom[13318] = 8'hf2 ;
            rom[13319] = 8'h0c ;
            rom[13320] = 8'hf7 ;
            rom[13321] = 8'h06 ;
            rom[13322] = 8'hf7 ;
            rom[13323] = 8'hfa ;
            rom[13324] = 8'h0b ;
            rom[13325] = 8'h2a ;
            rom[13326] = 8'hfb ;
            rom[13327] = 8'hf8 ;
            rom[13328] = 8'h08 ;
            rom[13329] = 8'hfb ;
            rom[13330] = 8'hff ;
            rom[13331] = 8'hfe ;
            rom[13332] = 8'h0a ;
            rom[13333] = 8'h03 ;
            rom[13334] = 8'h14 ;
            rom[13335] = 8'he5 ;
            rom[13336] = 8'h04 ;
            rom[13337] = 8'h07 ;
            rom[13338] = 8'h00 ;
            rom[13339] = 8'h26 ;
            rom[13340] = 8'he3 ;
            rom[13341] = 8'hef ;
            rom[13342] = 8'hf7 ;
            rom[13343] = 8'h14 ;
            rom[13344] = 8'hda ;
            rom[13345] = 8'hff ;
            rom[13346] = 8'h00 ;
            rom[13347] = 8'h13 ;
            rom[13348] = 8'hf8 ;
            rom[13349] = 8'h01 ;
            rom[13350] = 8'hcf ;
            rom[13351] = 8'hd5 ;
            rom[13352] = 8'hff ;
            rom[13353] = 8'h0d ;
            rom[13354] = 8'h06 ;
            rom[13355] = 8'he7 ;
            rom[13356] = 8'hfb ;
            rom[13357] = 8'h01 ;
            rom[13358] = 8'h02 ;
            rom[13359] = 8'h20 ;
            rom[13360] = 8'he1 ;
            rom[13361] = 8'h07 ;
            rom[13362] = 8'hfb ;
            rom[13363] = 8'he1 ;
            rom[13364] = 8'h00 ;
            rom[13365] = 8'hf8 ;
            rom[13366] = 8'h04 ;
            rom[13367] = 8'h06 ;
            rom[13368] = 8'h13 ;
            rom[13369] = 8'h1c ;
            rom[13370] = 8'hef ;
            rom[13371] = 8'hf5 ;
            rom[13372] = 8'hdf ;
            rom[13373] = 8'h08 ;
            rom[13374] = 8'h08 ;
            rom[13375] = 8'h16 ;
            rom[13376] = 8'h10 ;
            rom[13377] = 8'h00 ;
            rom[13378] = 8'h16 ;
            rom[13379] = 8'h06 ;
            rom[13380] = 8'h0f ;
            rom[13381] = 8'hfc ;
            rom[13382] = 8'h0b ;
            rom[13383] = 8'h30 ;
            rom[13384] = 8'hf8 ;
            rom[13385] = 8'h02 ;
            rom[13386] = 8'h0d ;
            rom[13387] = 8'hed ;
            rom[13388] = 8'hda ;
            rom[13389] = 8'hf0 ;
            rom[13390] = 8'h10 ;
            rom[13391] = 8'h07 ;
            rom[13392] = 8'hef ;
            rom[13393] = 8'he6 ;
            rom[13394] = 8'hee ;
            rom[13395] = 8'h07 ;
            rom[13396] = 8'hf3 ;
            rom[13397] = 8'hff ;
            rom[13398] = 8'h09 ;
            rom[13399] = 8'hde ;
            rom[13400] = 8'hfb ;
            rom[13401] = 8'hf0 ;
            rom[13402] = 8'he4 ;
            rom[13403] = 8'hec ;
            rom[13404] = 8'hfe ;
            rom[13405] = 8'h24 ;
            rom[13406] = 8'hfc ;
            rom[13407] = 8'h03 ;
            rom[13408] = 8'hf4 ;
            rom[13409] = 8'h08 ;
            rom[13410] = 8'hed ;
            rom[13411] = 8'hf1 ;
            rom[13412] = 8'h14 ;
            rom[13413] = 8'h00 ;
            rom[13414] = 8'h2b ;
            rom[13415] = 8'hdf ;
            rom[13416] = 8'h22 ;
            rom[13417] = 8'h05 ;
            rom[13418] = 8'hed ;
            rom[13419] = 8'h04 ;
            rom[13420] = 8'hd9 ;
            rom[13421] = 8'h0c ;
            rom[13422] = 8'h04 ;
            rom[13423] = 8'h16 ;
            rom[13424] = 8'h25 ;
            rom[13425] = 8'he7 ;
            rom[13426] = 8'h06 ;
            rom[13427] = 8'hf3 ;
            rom[13428] = 8'h2a ;
            rom[13429] = 8'hff ;
            rom[13430] = 8'hef ;
            rom[13431] = 8'h27 ;
            rom[13432] = 8'hd9 ;
            rom[13433] = 8'hdb ;
            rom[13434] = 8'h14 ;
            rom[13435] = 8'hf7 ;
            rom[13436] = 8'h1f ;
            rom[13437] = 8'he0 ;
            rom[13438] = 8'heb ;
            rom[13439] = 8'h07 ;
            rom[13440] = 8'h09 ;
            rom[13441] = 8'hfd ;
            rom[13442] = 8'hfa ;
            rom[13443] = 8'hfc ;
            rom[13444] = 8'h02 ;
            rom[13445] = 8'hfc ;
            rom[13446] = 8'hed ;
            rom[13447] = 8'h09 ;
            rom[13448] = 8'he6 ;
            rom[13449] = 8'hf5 ;
            rom[13450] = 8'h0e ;
            rom[13451] = 8'h11 ;
            rom[13452] = 8'he6 ;
            rom[13453] = 8'h06 ;
            rom[13454] = 8'hf6 ;
            rom[13455] = 8'hfb ;
            rom[13456] = 8'h0d ;
            rom[13457] = 8'h07 ;
            rom[13458] = 8'h28 ;
            rom[13459] = 8'h18 ;
            rom[13460] = 8'hf0 ;
            rom[13461] = 8'he9 ;
            rom[13462] = 8'hf9 ;
            rom[13463] = 8'hfe ;
            rom[13464] = 8'h01 ;
            rom[13465] = 8'hff ;
            rom[13466] = 8'h0b ;
            rom[13467] = 8'h00 ;
            rom[13468] = 8'hcc ;
            rom[13469] = 8'hfe ;
            rom[13470] = 8'h22 ;
            rom[13471] = 8'h0c ;
            rom[13472] = 8'hbe ;
            rom[13473] = 8'h11 ;
            rom[13474] = 8'hfa ;
            rom[13475] = 8'h01 ;
            rom[13476] = 8'h1d ;
            rom[13477] = 8'h12 ;
            rom[13478] = 8'hff ;
            rom[13479] = 8'h26 ;
            rom[13480] = 8'h11 ;
            rom[13481] = 8'h06 ;
            rom[13482] = 8'h02 ;
            rom[13483] = 8'hf2 ;
            rom[13484] = 8'hda ;
            rom[13485] = 8'hfa ;
            rom[13486] = 8'h13 ;
            rom[13487] = 8'hd2 ;
            rom[13488] = 8'h0c ;
            rom[13489] = 8'h14 ;
            rom[13490] = 8'he1 ;
            rom[13491] = 8'h22 ;
            rom[13492] = 8'he7 ;
            rom[13493] = 8'h0a ;
            rom[13494] = 8'h01 ;
            rom[13495] = 8'h0c ;
            rom[13496] = 8'he9 ;
            rom[13497] = 8'h17 ;
            rom[13498] = 8'hf6 ;
            rom[13499] = 8'h08 ;
            rom[13500] = 8'hc5 ;
            rom[13501] = 8'he9 ;
            rom[13502] = 8'he6 ;
            rom[13503] = 8'h13 ;
            rom[13504] = 8'h01 ;
            rom[13505] = 8'hee ;
            rom[13506] = 8'hff ;
            rom[13507] = 8'h12 ;
            rom[13508] = 8'he2 ;
            rom[13509] = 8'hfb ;
            rom[13510] = 8'h0c ;
            rom[13511] = 8'h10 ;
            rom[13512] = 8'h0f ;
            rom[13513] = 8'h10 ;
            rom[13514] = 8'hf3 ;
            rom[13515] = 8'hfd ;
            rom[13516] = 8'hd4 ;
            rom[13517] = 8'h13 ;
            rom[13518] = 8'h05 ;
            rom[13519] = 8'h00 ;
            rom[13520] = 8'hdb ;
            rom[13521] = 8'hf3 ;
            rom[13522] = 8'h04 ;
            rom[13523] = 8'hfc ;
            rom[13524] = 8'hf1 ;
            rom[13525] = 8'h0f ;
            rom[13526] = 8'hf9 ;
            rom[13527] = 8'hfa ;
            rom[13528] = 8'h0d ;
            rom[13529] = 8'hf5 ;
            rom[13530] = 8'hed ;
            rom[13531] = 8'h2f ;
            rom[13532] = 8'hcc ;
            rom[13533] = 8'h02 ;
            rom[13534] = 8'h0f ;
            rom[13535] = 8'h10 ;
            rom[13536] = 8'hea ;
            rom[13537] = 8'hfc ;
            rom[13538] = 8'h0d ;
            rom[13539] = 8'h08 ;
            rom[13540] = 8'hf6 ;
            rom[13541] = 8'h04 ;
            rom[13542] = 8'h10 ;
            rom[13543] = 8'hf4 ;
            rom[13544] = 8'h0f ;
            rom[13545] = 8'hfd ;
            rom[13546] = 8'hb1 ;
            rom[13547] = 8'h11 ;
            rom[13548] = 8'hf4 ;
            rom[13549] = 8'hf9 ;
            rom[13550] = 8'heb ;
            rom[13551] = 8'h0d ;
            rom[13552] = 8'h1f ;
            rom[13553] = 8'hf4 ;
            rom[13554] = 8'h22 ;
            rom[13555] = 8'hfe ;
            rom[13556] = 8'h06 ;
            rom[13557] = 8'hff ;
            rom[13558] = 8'hc0 ;
            rom[13559] = 8'h19 ;
            rom[13560] = 8'hfb ;
            rom[13561] = 8'hf4 ;
            rom[13562] = 8'hff ;
            rom[13563] = 8'h08 ;
            rom[13564] = 8'h1e ;
            rom[13565] = 8'h09 ;
            rom[13566] = 8'h08 ;
            rom[13567] = 8'hf8 ;
            rom[13568] = 8'h10 ;
            rom[13569] = 8'hf5 ;
            rom[13570] = 8'h0b ;
            rom[13571] = 8'hf3 ;
            rom[13572] = 8'h04 ;
            rom[13573] = 8'h11 ;
            rom[13574] = 8'hfa ;
            rom[13575] = 8'h02 ;
            rom[13576] = 8'hfd ;
            rom[13577] = 8'h11 ;
            rom[13578] = 8'h13 ;
            rom[13579] = 8'hfb ;
            rom[13580] = 8'h09 ;
            rom[13581] = 8'h39 ;
            rom[13582] = 8'hc9 ;
            rom[13583] = 8'hf4 ;
            rom[13584] = 8'h07 ;
            rom[13585] = 8'hff ;
            rom[13586] = 8'hf4 ;
            rom[13587] = 8'h0b ;
            rom[13588] = 8'h0c ;
            rom[13589] = 8'hdb ;
            rom[13590] = 8'hf3 ;
            rom[13591] = 8'hff ;
            rom[13592] = 8'hf5 ;
            rom[13593] = 8'hd3 ;
            rom[13594] = 8'hf2 ;
            rom[13595] = 8'h0c ;
            rom[13596] = 8'hf7 ;
            rom[13597] = 8'h03 ;
            rom[13598] = 8'h05 ;
            rom[13599] = 8'h13 ;
            rom[13600] = 8'hd5 ;
            rom[13601] = 8'h12 ;
            rom[13602] = 8'h19 ;
            rom[13603] = 8'hf6 ;
            rom[13604] = 8'h0e ;
            rom[13605] = 8'h0b ;
            rom[13606] = 8'hd9 ;
            rom[13607] = 8'he2 ;
            rom[13608] = 8'h10 ;
            rom[13609] = 8'hf6 ;
            rom[13610] = 8'hed ;
            rom[13611] = 8'h0e ;
            rom[13612] = 8'h03 ;
            rom[13613] = 8'h04 ;
            rom[13614] = 8'hfe ;
            rom[13615] = 8'h04 ;
            rom[13616] = 8'he4 ;
            rom[13617] = 8'hf1 ;
            rom[13618] = 8'hf9 ;
            rom[13619] = 8'hf6 ;
            rom[13620] = 8'hf9 ;
            rom[13621] = 8'he9 ;
            rom[13622] = 8'h0b ;
            rom[13623] = 8'h09 ;
            rom[13624] = 8'h10 ;
            rom[13625] = 8'h04 ;
            rom[13626] = 8'hdd ;
            rom[13627] = 8'he9 ;
            rom[13628] = 8'h02 ;
            rom[13629] = 8'hee ;
            rom[13630] = 8'h11 ;
            rom[13631] = 8'heb ;
            rom[13632] = 8'h17 ;
            rom[13633] = 8'h03 ;
            rom[13634] = 8'h01 ;
            rom[13635] = 8'h12 ;
            rom[13636] = 8'h0e ;
            rom[13637] = 8'hf1 ;
            rom[13638] = 8'hf9 ;
            rom[13639] = 8'h13 ;
            rom[13640] = 8'hfb ;
            rom[13641] = 8'hfc ;
            rom[13642] = 8'hf4 ;
            rom[13643] = 8'hd6 ;
            rom[13644] = 8'hf4 ;
            rom[13645] = 8'h01 ;
            rom[13646] = 8'hfb ;
            rom[13647] = 8'hca ;
            rom[13648] = 8'hd7 ;
            rom[13649] = 8'h04 ;
            rom[13650] = 8'h13 ;
            rom[13651] = 8'h0d ;
            rom[13652] = 8'h03 ;
            rom[13653] = 8'hfd ;
            rom[13654] = 8'h2b ;
            rom[13655] = 8'h19 ;
            rom[13656] = 8'hf8 ;
            rom[13657] = 8'h12 ;
            rom[13658] = 8'h16 ;
            rom[13659] = 8'h02 ;
            rom[13660] = 8'hea ;
            rom[13661] = 8'hef ;
            rom[13662] = 8'hf9 ;
            rom[13663] = 8'h12 ;
            rom[13664] = 8'hdc ;
            rom[13665] = 8'hfd ;
            rom[13666] = 8'hd8 ;
            rom[13667] = 8'h19 ;
            rom[13668] = 8'h09 ;
            rom[13669] = 8'h01 ;
            rom[13670] = 8'h00 ;
            rom[13671] = 8'he0 ;
            rom[13672] = 8'hf0 ;
            rom[13673] = 8'h1c ;
            rom[13674] = 8'h1e ;
            rom[13675] = 8'h02 ;
            rom[13676] = 8'hf2 ;
            rom[13677] = 8'h13 ;
            rom[13678] = 8'hfc ;
            rom[13679] = 8'h29 ;
            rom[13680] = 8'hf1 ;
            rom[13681] = 8'h26 ;
            rom[13682] = 8'h01 ;
            rom[13683] = 8'hfb ;
            rom[13684] = 8'hf4 ;
            rom[13685] = 8'h16 ;
            rom[13686] = 8'hfe ;
            rom[13687] = 8'h15 ;
            rom[13688] = 8'hf7 ;
            rom[13689] = 8'hfb ;
            rom[13690] = 8'h05 ;
            rom[13691] = 8'hec ;
            rom[13692] = 8'h08 ;
            rom[13693] = 8'h10 ;
            rom[13694] = 8'h1e ;
            rom[13695] = 8'h1a ;
            rom[13696] = 8'h06 ;
            rom[13697] = 8'h01 ;
            rom[13698] = 8'h00 ;
            rom[13699] = 8'h12 ;
            rom[13700] = 8'hf7 ;
            rom[13701] = 8'h0b ;
            rom[13702] = 8'h05 ;
            rom[13703] = 8'h0e ;
            rom[13704] = 8'hf9 ;
            rom[13705] = 8'hf9 ;
            rom[13706] = 8'h00 ;
            rom[13707] = 8'hf6 ;
            rom[13708] = 8'h00 ;
            rom[13709] = 8'h09 ;
            rom[13710] = 8'h04 ;
            rom[13711] = 8'hc5 ;
            rom[13712] = 8'hcd ;
            rom[13713] = 8'h03 ;
            rom[13714] = 8'hfb ;
            rom[13715] = 8'hf1 ;
            rom[13716] = 8'hfa ;
            rom[13717] = 8'he0 ;
            rom[13718] = 8'hd7 ;
            rom[13719] = 8'h19 ;
            rom[13720] = 8'h14 ;
            rom[13721] = 8'he1 ;
            rom[13722] = 8'hdf ;
            rom[13723] = 8'h19 ;
            rom[13724] = 8'h04 ;
            rom[13725] = 8'h00 ;
            rom[13726] = 8'h02 ;
            rom[13727] = 8'hfb ;
            rom[13728] = 8'h06 ;
            rom[13729] = 8'hf9 ;
            rom[13730] = 8'hd6 ;
            rom[13731] = 8'h02 ;
            rom[13732] = 8'h02 ;
            rom[13733] = 8'hf8 ;
            rom[13734] = 8'h12 ;
            rom[13735] = 8'h1e ;
            rom[13736] = 8'hfc ;
            rom[13737] = 8'hee ;
            rom[13738] = 8'hf7 ;
            rom[13739] = 8'h2a ;
            rom[13740] = 8'hef ;
            rom[13741] = 8'h01 ;
            rom[13742] = 8'h0d ;
            rom[13743] = 8'hc5 ;
            rom[13744] = 8'hd7 ;
            rom[13745] = 8'hf8 ;
            rom[13746] = 8'h0c ;
            rom[13747] = 8'hfe ;
            rom[13748] = 8'hdf ;
            rom[13749] = 8'hf4 ;
            rom[13750] = 8'h14 ;
            rom[13751] = 8'h14 ;
            rom[13752] = 8'h0d ;
            rom[13753] = 8'hf6 ;
            rom[13754] = 8'h0e ;
            rom[13755] = 8'h07 ;
            rom[13756] = 8'h0f ;
            rom[13757] = 8'hcc ;
            rom[13758] = 8'h0a ;
            rom[13759] = 8'hf7 ;
            rom[13760] = 8'hf6 ;
            rom[13761] = 8'h10 ;
            rom[13762] = 8'h04 ;
            rom[13763] = 8'hfc ;
            rom[13764] = 8'h0b ;
            rom[13765] = 8'h0f ;
            rom[13766] = 8'h14 ;
            rom[13767] = 8'h20 ;
            rom[13768] = 8'h0c ;
            rom[13769] = 8'h1f ;
            rom[13770] = 8'hf5 ;
            rom[13771] = 8'he7 ;
            rom[13772] = 8'hf8 ;
            rom[13773] = 8'h0a ;
            rom[13774] = 8'hfb ;
            rom[13775] = 8'he3 ;
            rom[13776] = 8'hea ;
            rom[13777] = 8'hfa ;
            rom[13778] = 8'h22 ;
            rom[13779] = 8'h15 ;
            rom[13780] = 8'h1b ;
            rom[13781] = 8'hfc ;
            rom[13782] = 8'hf6 ;
            rom[13783] = 8'h13 ;
            rom[13784] = 8'h18 ;
            rom[13785] = 8'h18 ;
            rom[13786] = 8'h23 ;
            rom[13787] = 8'heb ;
            rom[13788] = 8'hd1 ;
            rom[13789] = 8'hfe ;
            rom[13790] = 8'hfe ;
            rom[13791] = 8'h04 ;
            rom[13792] = 8'he2 ;
            rom[13793] = 8'hff ;
            rom[13794] = 8'h1b ;
            rom[13795] = 8'hf9 ;
            rom[13796] = 8'h0c ;
            rom[13797] = 8'he2 ;
            rom[13798] = 8'hfe ;
            rom[13799] = 8'hdf ;
            rom[13800] = 8'h0c ;
            rom[13801] = 8'h03 ;
            rom[13802] = 8'h14 ;
            rom[13803] = 8'h1b ;
            rom[13804] = 8'h00 ;
            rom[13805] = 8'h0f ;
            rom[13806] = 8'h21 ;
            rom[13807] = 8'h36 ;
            rom[13808] = 8'hfc ;
            rom[13809] = 8'h14 ;
            rom[13810] = 8'h15 ;
            rom[13811] = 8'h0e ;
            rom[13812] = 8'hee ;
            rom[13813] = 8'h09 ;
            rom[13814] = 8'h17 ;
            rom[13815] = 8'h17 ;
            rom[13816] = 8'he5 ;
            rom[13817] = 8'hfb ;
            rom[13818] = 8'h0c ;
            rom[13819] = 8'h0d ;
            rom[13820] = 8'h03 ;
            rom[13821] = 8'h06 ;
            rom[13822] = 8'hf5 ;
            rom[13823] = 8'h03 ;
            rom[13824] = 8'h1a ;
            rom[13825] = 8'hf0 ;
            rom[13826] = 8'h18 ;
            rom[13827] = 8'h09 ;
            rom[13828] = 8'hea ;
            rom[13829] = 8'h07 ;
            rom[13830] = 8'hf6 ;
            rom[13831] = 8'hfa ;
            rom[13832] = 8'hcf ;
            rom[13833] = 8'h0e ;
            rom[13834] = 8'h13 ;
            rom[13835] = 8'hfd ;
            rom[13836] = 8'h05 ;
            rom[13837] = 8'h0d ;
            rom[13838] = 8'hdd ;
            rom[13839] = 8'hc9 ;
            rom[13840] = 8'hd5 ;
            rom[13841] = 8'h03 ;
            rom[13842] = 8'hf1 ;
            rom[13843] = 8'h12 ;
            rom[13844] = 8'hfe ;
            rom[13845] = 8'h07 ;
            rom[13846] = 8'hfa ;
            rom[13847] = 8'h13 ;
            rom[13848] = 8'h0b ;
            rom[13849] = 8'hcd ;
            rom[13850] = 8'hdd ;
            rom[13851] = 8'hfa ;
            rom[13852] = 8'hec ;
            rom[13853] = 8'hf1 ;
            rom[13854] = 8'h0b ;
            rom[13855] = 8'hf6 ;
            rom[13856] = 8'hd5 ;
            rom[13857] = 8'hf0 ;
            rom[13858] = 8'hd0 ;
            rom[13859] = 8'h0d ;
            rom[13860] = 8'hfb ;
            rom[13861] = 8'hf9 ;
            rom[13862] = 8'h13 ;
            rom[13863] = 8'h04 ;
            rom[13864] = 8'h18 ;
            rom[13865] = 8'hf3 ;
            rom[13866] = 8'h0c ;
            rom[13867] = 8'h17 ;
            rom[13868] = 8'hf4 ;
            rom[13869] = 8'hfa ;
            rom[13870] = 8'h19 ;
            rom[13871] = 8'hf7 ;
            rom[13872] = 8'h08 ;
            rom[13873] = 8'hec ;
            rom[13874] = 8'h06 ;
            rom[13875] = 8'hf1 ;
            rom[13876] = 8'h01 ;
            rom[13877] = 8'h08 ;
            rom[13878] = 8'hf7 ;
            rom[13879] = 8'h20 ;
            rom[13880] = 8'hff ;
            rom[13881] = 8'hd2 ;
            rom[13882] = 8'h07 ;
            rom[13883] = 8'h0f ;
            rom[13884] = 8'hfc ;
            rom[13885] = 8'he8 ;
            rom[13886] = 8'h08 ;
            rom[13887] = 8'h12 ;
            rom[13888] = 8'h04 ;
            rom[13889] = 8'h01 ;
            rom[13890] = 8'h00 ;
            rom[13891] = 8'h25 ;
            rom[13892] = 8'hd5 ;
            rom[13893] = 8'hff ;
            rom[13894] = 8'h02 ;
            rom[13895] = 8'hff ;
            rom[13896] = 8'he8 ;
            rom[13897] = 8'h01 ;
            rom[13898] = 8'h14 ;
            rom[13899] = 8'h04 ;
            rom[13900] = 8'hf6 ;
            rom[13901] = 8'h0d ;
            rom[13902] = 8'hf2 ;
            rom[13903] = 8'hdd ;
            rom[13904] = 8'hb0 ;
            rom[13905] = 8'h05 ;
            rom[13906] = 8'h07 ;
            rom[13907] = 8'hf3 ;
            rom[13908] = 8'hf7 ;
            rom[13909] = 8'h17 ;
            rom[13910] = 8'hf0 ;
            rom[13911] = 8'hf1 ;
            rom[13912] = 8'h08 ;
            rom[13913] = 8'hd6 ;
            rom[13914] = 8'hf4 ;
            rom[13915] = 8'h1e ;
            rom[13916] = 8'hde ;
            rom[13917] = 8'h24 ;
            rom[13918] = 8'h06 ;
            rom[13919] = 8'hf4 ;
            rom[13920] = 8'h1b ;
            rom[13921] = 8'he4 ;
            rom[13922] = 8'h1e ;
            rom[13923] = 8'h09 ;
            rom[13924] = 8'h00 ;
            rom[13925] = 8'h03 ;
            rom[13926] = 8'h10 ;
            rom[13927] = 8'hf1 ;
            rom[13928] = 8'h03 ;
            rom[13929] = 8'hc9 ;
            rom[13930] = 8'hc8 ;
            rom[13931] = 8'h25 ;
            rom[13932] = 8'h03 ;
            rom[13933] = 8'hf6 ;
            rom[13934] = 8'h00 ;
            rom[13935] = 8'h01 ;
            rom[13936] = 8'h0a ;
            rom[13937] = 8'hfd ;
            rom[13938] = 8'h15 ;
            rom[13939] = 8'hf5 ;
            rom[13940] = 8'hfe ;
            rom[13941] = 8'h06 ;
            rom[13942] = 8'hd6 ;
            rom[13943] = 8'h05 ;
            rom[13944] = 8'h0c ;
            rom[13945] = 8'hf2 ;
            rom[13946] = 8'h0c ;
            rom[13947] = 8'h14 ;
            rom[13948] = 8'h19 ;
            rom[13949] = 8'hff ;
            rom[13950] = 8'h1c ;
            rom[13951] = 8'hfc ;
            rom[13952] = 8'h09 ;
            rom[13953] = 8'h14 ;
            rom[13954] = 8'he6 ;
            rom[13955] = 8'h1c ;
            rom[13956] = 8'hff ;
            rom[13957] = 8'hf7 ;
            rom[13958] = 8'h04 ;
            rom[13959] = 8'h07 ;
            rom[13960] = 8'hf9 ;
            rom[13961] = 8'he6 ;
            rom[13962] = 8'h06 ;
            rom[13963] = 8'hec ;
            rom[13964] = 8'h1f ;
            rom[13965] = 8'h0f ;
            rom[13966] = 8'h05 ;
            rom[13967] = 8'heb ;
            rom[13968] = 8'hb9 ;
            rom[13969] = 8'h03 ;
            rom[13970] = 8'h13 ;
            rom[13971] = 8'hde ;
            rom[13972] = 8'h02 ;
            rom[13973] = 8'hed ;
            rom[13974] = 8'h1d ;
            rom[13975] = 8'h0c ;
            rom[13976] = 8'h00 ;
            rom[13977] = 8'hfb ;
            rom[13978] = 8'h00 ;
            rom[13979] = 8'h18 ;
            rom[13980] = 8'hf5 ;
            rom[13981] = 8'hfd ;
            rom[13982] = 8'hf1 ;
            rom[13983] = 8'h18 ;
            rom[13984] = 8'h0e ;
            rom[13985] = 8'hf5 ;
            rom[13986] = 8'hfd ;
            rom[13987] = 8'hd3 ;
            rom[13988] = 8'h12 ;
            rom[13989] = 8'hff ;
            rom[13990] = 8'h11 ;
            rom[13991] = 8'hf9 ;
            rom[13992] = 8'h10 ;
            rom[13993] = 8'hde ;
            rom[13994] = 8'h02 ;
            rom[13995] = 8'h19 ;
            rom[13996] = 8'hff ;
            rom[13997] = 8'hfd ;
            rom[13998] = 8'hff ;
            rom[13999] = 8'h00 ;
            rom[14000] = 8'h02 ;
            rom[14001] = 8'h05 ;
            rom[14002] = 8'h11 ;
            rom[14003] = 8'hfa ;
            rom[14004] = 8'hff ;
            rom[14005] = 8'h05 ;
            rom[14006] = 8'h00 ;
            rom[14007] = 8'hff ;
            rom[14008] = 8'h09 ;
            rom[14009] = 8'h0f ;
            rom[14010] = 8'h18 ;
            rom[14011] = 8'h03 ;
            rom[14012] = 8'h0d ;
            rom[14013] = 8'h23 ;
            rom[14014] = 8'h05 ;
            rom[14015] = 8'h06 ;
            rom[14016] = 8'he5 ;
            rom[14017] = 8'h0f ;
            rom[14018] = 8'h0b ;
            rom[14019] = 8'h08 ;
            rom[14020] = 8'hf0 ;
            rom[14021] = 8'he0 ;
            rom[14022] = 8'h0e ;
            rom[14023] = 8'hfd ;
            rom[14024] = 8'h01 ;
            rom[14025] = 8'h09 ;
            rom[14026] = 8'he7 ;
            rom[14027] = 8'h08 ;
            rom[14028] = 8'h0c ;
            rom[14029] = 8'h04 ;
            rom[14030] = 8'h0a ;
            rom[14031] = 8'hd7 ;
            rom[14032] = 8'hd4 ;
            rom[14033] = 8'hf8 ;
            rom[14034] = 8'hf5 ;
            rom[14035] = 8'h05 ;
            rom[14036] = 8'h10 ;
            rom[14037] = 8'hcf ;
            rom[14038] = 8'he9 ;
            rom[14039] = 8'h10 ;
            rom[14040] = 8'hfc ;
            rom[14041] = 8'hea ;
            rom[14042] = 8'hf6 ;
            rom[14043] = 8'hfe ;
            rom[14044] = 8'hca ;
            rom[14045] = 8'hfe ;
            rom[14046] = 8'h0a ;
            rom[14047] = 8'h0f ;
            rom[14048] = 8'h01 ;
            rom[14049] = 8'h08 ;
            rom[14050] = 8'h16 ;
            rom[14051] = 8'hfe ;
            rom[14052] = 8'h20 ;
            rom[14053] = 8'hfa ;
            rom[14054] = 8'h1d ;
            rom[14055] = 8'hf1 ;
            rom[14056] = 8'h14 ;
            rom[14057] = 8'hfd ;
            rom[14058] = 8'hfc ;
            rom[14059] = 8'h07 ;
            rom[14060] = 8'h0a ;
            rom[14061] = 8'h01 ;
            rom[14062] = 8'hf0 ;
            rom[14063] = 8'h01 ;
            rom[14064] = 8'h19 ;
            rom[14065] = 8'h08 ;
            rom[14066] = 8'heb ;
            rom[14067] = 8'hfa ;
            rom[14068] = 8'hfc ;
            rom[14069] = 8'hf3 ;
            rom[14070] = 8'h0d ;
            rom[14071] = 8'h20 ;
            rom[14072] = 8'hfe ;
            rom[14073] = 8'heb ;
            rom[14074] = 8'heb ;
            rom[14075] = 8'h02 ;
            rom[14076] = 8'h10 ;
            rom[14077] = 8'h03 ;
            rom[14078] = 8'h10 ;
            rom[14079] = 8'h0c ;
            rom[14080] = 8'hfc ;
            rom[14081] = 8'h02 ;
            rom[14082] = 8'hfe ;
            rom[14083] = 8'h14 ;
            rom[14084] = 8'h01 ;
            rom[14085] = 8'h1b ;
            rom[14086] = 8'h09 ;
            rom[14087] = 8'h19 ;
            rom[14088] = 8'he2 ;
            rom[14089] = 8'h19 ;
            rom[14090] = 8'hf9 ;
            rom[14091] = 8'hef ;
            rom[14092] = 8'h0c ;
            rom[14093] = 8'h17 ;
            rom[14094] = 8'hf6 ;
            rom[14095] = 8'hec ;
            rom[14096] = 8'hf6 ;
            rom[14097] = 8'h1e ;
            rom[14098] = 8'h04 ;
            rom[14099] = 8'h1d ;
            rom[14100] = 8'h10 ;
            rom[14101] = 8'hf3 ;
            rom[14102] = 8'h0e ;
            rom[14103] = 8'h14 ;
            rom[14104] = 8'h07 ;
            rom[14105] = 8'hf7 ;
            rom[14106] = 8'h13 ;
            rom[14107] = 8'h08 ;
            rom[14108] = 8'h17 ;
            rom[14109] = 8'hd7 ;
            rom[14110] = 8'hf6 ;
            rom[14111] = 8'h16 ;
            rom[14112] = 8'hc3 ;
            rom[14113] = 8'h04 ;
            rom[14114] = 8'h16 ;
            rom[14115] = 8'h1d ;
            rom[14116] = 8'h12 ;
            rom[14117] = 8'hf3 ;
            rom[14118] = 8'heb ;
            rom[14119] = 8'hf9 ;
            rom[14120] = 8'hf8 ;
            rom[14121] = 8'h04 ;
            rom[14122] = 8'h02 ;
            rom[14123] = 8'h09 ;
            rom[14124] = 8'hfa ;
            rom[14125] = 8'h23 ;
            rom[14126] = 8'hfa ;
            rom[14127] = 8'h28 ;
            rom[14128] = 8'heb ;
            rom[14129] = 8'h1c ;
            rom[14130] = 8'hfc ;
            rom[14131] = 8'h05 ;
            rom[14132] = 8'h00 ;
            rom[14133] = 8'he6 ;
            rom[14134] = 8'h11 ;
            rom[14135] = 8'h1a ;
            rom[14136] = 8'hfe ;
            rom[14137] = 8'hff ;
            rom[14138] = 8'h02 ;
            rom[14139] = 8'hff ;
            rom[14140] = 8'h00 ;
            rom[14141] = 8'hff ;
            rom[14142] = 8'hfc ;
            rom[14143] = 8'h15 ;
            rom[14144] = 8'h18 ;
            rom[14145] = 8'h05 ;
            rom[14146] = 8'h01 ;
            rom[14147] = 8'hed ;
            rom[14148] = 8'h13 ;
            rom[14149] = 8'h09 ;
            rom[14150] = 8'h11 ;
            rom[14151] = 8'he9 ;
            rom[14152] = 8'h10 ;
            rom[14153] = 8'hf2 ;
            rom[14154] = 8'h0f ;
            rom[14155] = 8'h02 ;
            rom[14156] = 8'he1 ;
            rom[14157] = 8'h16 ;
            rom[14158] = 8'h0b ;
            rom[14159] = 8'hec ;
            rom[14160] = 8'h10 ;
            rom[14161] = 8'h2f ;
            rom[14162] = 8'he4 ;
            rom[14163] = 8'hf6 ;
            rom[14164] = 8'hd4 ;
            rom[14165] = 8'he1 ;
            rom[14166] = 8'hfb ;
            rom[14167] = 8'hff ;
            rom[14168] = 8'hf7 ;
            rom[14169] = 8'h02 ;
            rom[14170] = 8'h0d ;
            rom[14171] = 8'h0a ;
            rom[14172] = 8'h1b ;
            rom[14173] = 8'hf4 ;
            rom[14174] = 8'h02 ;
            rom[14175] = 8'h08 ;
            rom[14176] = 8'hf4 ;
            rom[14177] = 8'h16 ;
            rom[14178] = 8'h05 ;
            rom[14179] = 8'hf2 ;
            rom[14180] = 8'h11 ;
            rom[14181] = 8'hfc ;
            rom[14182] = 8'hf2 ;
            rom[14183] = 8'hd0 ;
            rom[14184] = 8'h18 ;
            rom[14185] = 8'hfa ;
            rom[14186] = 8'h0b ;
            rom[14187] = 8'h0e ;
            rom[14188] = 8'hef ;
            rom[14189] = 8'hfc ;
            rom[14190] = 8'heb ;
            rom[14191] = 8'h04 ;
            rom[14192] = 8'h06 ;
            rom[14193] = 8'hd1 ;
            rom[14194] = 8'h03 ;
            rom[14195] = 8'hda ;
            rom[14196] = 8'h01 ;
            rom[14197] = 8'hf6 ;
            rom[14198] = 8'hea ;
            rom[14199] = 8'h1b ;
            rom[14200] = 8'hf6 ;
            rom[14201] = 8'h05 ;
            rom[14202] = 8'h08 ;
            rom[14203] = 8'hf5 ;
            rom[14204] = 8'h14 ;
            rom[14205] = 8'hfb ;
            rom[14206] = 8'hee ;
            rom[14207] = 8'h19 ;
            rom[14208] = 8'h1b ;
            rom[14209] = 8'hfa ;
            rom[14210] = 8'hdb ;
            rom[14211] = 8'h12 ;
            rom[14212] = 8'hf0 ;
            rom[14213] = 8'hf9 ;
            rom[14214] = 8'hf2 ;
            rom[14215] = 8'hfa ;
            rom[14216] = 8'h00 ;
            rom[14217] = 8'h09 ;
            rom[14218] = 8'h07 ;
            rom[14219] = 8'h07 ;
            rom[14220] = 8'h14 ;
            rom[14221] = 8'h06 ;
            rom[14222] = 8'hf8 ;
            rom[14223] = 8'hee ;
            rom[14224] = 8'h02 ;
            rom[14225] = 8'hfb ;
            rom[14226] = 8'h10 ;
            rom[14227] = 8'hff ;
            rom[14228] = 8'h09 ;
            rom[14229] = 8'h01 ;
            rom[14230] = 8'hf4 ;
            rom[14231] = 8'h09 ;
            rom[14232] = 8'h0a ;
            rom[14233] = 8'h02 ;
            rom[14234] = 8'h30 ;
            rom[14235] = 8'h05 ;
            rom[14236] = 8'hf9 ;
            rom[14237] = 8'hde ;
            rom[14238] = 8'hf6 ;
            rom[14239] = 8'hd9 ;
            rom[14240] = 8'hd6 ;
            rom[14241] = 8'hf6 ;
            rom[14242] = 8'hfe ;
            rom[14243] = 8'h04 ;
            rom[14244] = 8'heb ;
            rom[14245] = 8'h13 ;
            rom[14246] = 8'he9 ;
            rom[14247] = 8'h0c ;
            rom[14248] = 8'h0e ;
            rom[14249] = 8'h02 ;
            rom[14250] = 8'h03 ;
            rom[14251] = 8'h07 ;
            rom[14252] = 8'heb ;
            rom[14253] = 8'h19 ;
            rom[14254] = 8'hfe ;
            rom[14255] = 8'he5 ;
            rom[14256] = 8'hf6 ;
            rom[14257] = 8'hf4 ;
            rom[14258] = 8'h02 ;
            rom[14259] = 8'h18 ;
            rom[14260] = 8'h0d ;
            rom[14261] = 8'h04 ;
            rom[14262] = 8'h15 ;
            rom[14263] = 8'h0b ;
            rom[14264] = 8'h0c ;
            rom[14265] = 8'h10 ;
            rom[14266] = 8'h2c ;
            rom[14267] = 8'h11 ;
            rom[14268] = 8'hfd ;
            rom[14269] = 8'hd9 ;
            rom[14270] = 8'h0c ;
            rom[14271] = 8'h07 ;
            rom[14272] = 8'he3 ;
            rom[14273] = 8'hf7 ;
            rom[14274] = 8'he7 ;
            rom[14275] = 8'h00 ;
            rom[14276] = 8'h11 ;
            rom[14277] = 8'h10 ;
            rom[14278] = 8'h00 ;
            rom[14279] = 8'h0e ;
            rom[14280] = 8'h1f ;
            rom[14281] = 8'hfa ;
            rom[14282] = 8'h11 ;
            rom[14283] = 8'h09 ;
            rom[14284] = 8'h07 ;
            rom[14285] = 8'he0 ;
            rom[14286] = 8'h0b ;
            rom[14287] = 8'hda ;
            rom[14288] = 8'hfa ;
            rom[14289] = 8'h24 ;
            rom[14290] = 8'hfb ;
            rom[14291] = 8'hfc ;
            rom[14292] = 8'heb ;
            rom[14293] = 8'hf5 ;
            rom[14294] = 8'h00 ;
            rom[14295] = 8'h0f ;
            rom[14296] = 8'hda ;
            rom[14297] = 8'h30 ;
            rom[14298] = 8'h12 ;
            rom[14299] = 8'h03 ;
            rom[14300] = 8'h08 ;
            rom[14301] = 8'he2 ;
            rom[14302] = 8'hce ;
            rom[14303] = 8'h17 ;
            rom[14304] = 8'h0d ;
            rom[14305] = 8'h16 ;
            rom[14306] = 8'hf7 ;
            rom[14307] = 8'hf5 ;
            rom[14308] = 8'h1a ;
            rom[14309] = 8'hee ;
            rom[14310] = 8'h09 ;
            rom[14311] = 8'he3 ;
            rom[14312] = 8'h05 ;
            rom[14313] = 8'h07 ;
            rom[14314] = 8'h1c ;
            rom[14315] = 8'h1b ;
            rom[14316] = 8'hf9 ;
            rom[14317] = 8'h07 ;
            rom[14318] = 8'h0b ;
            rom[14319] = 8'h18 ;
            rom[14320] = 8'h07 ;
            rom[14321] = 8'hf5 ;
            rom[14322] = 8'h07 ;
            rom[14323] = 8'hc3 ;
            rom[14324] = 8'he5 ;
            rom[14325] = 8'h1e ;
            rom[14326] = 8'h05 ;
            rom[14327] = 8'h02 ;
            rom[14328] = 8'hff ;
            rom[14329] = 8'h07 ;
            rom[14330] = 8'h12 ;
            rom[14331] = 8'hf3 ;
            rom[14332] = 8'h0f ;
            rom[14333] = 8'h1b ;
            rom[14334] = 8'hea ;
            rom[14335] = 8'h01 ;
            rom[14336] = 8'h17 ;
            rom[14337] = 8'hf9 ;
            rom[14338] = 8'hf0 ;
            rom[14339] = 8'he5 ;
            rom[14340] = 8'h17 ;
            rom[14341] = 8'h0f ;
            rom[14342] = 8'h20 ;
            rom[14343] = 8'hcf ;
            rom[14344] = 8'hfe ;
            rom[14345] = 8'h01 ;
            rom[14346] = 8'he0 ;
            rom[14347] = 8'h08 ;
            rom[14348] = 8'hd3 ;
            rom[14349] = 8'hf9 ;
            rom[14350] = 8'h00 ;
            rom[14351] = 8'hf4 ;
            rom[14352] = 8'h02 ;
            rom[14353] = 8'h0f ;
            rom[14354] = 8'hfe ;
            rom[14355] = 8'h05 ;
            rom[14356] = 8'hfd ;
            rom[14357] = 8'h0a ;
            rom[14358] = 8'hd9 ;
            rom[14359] = 8'hf2 ;
            rom[14360] = 8'hf7 ;
            rom[14361] = 8'he6 ;
            rom[14362] = 8'hf7 ;
            rom[14363] = 8'he8 ;
            rom[14364] = 8'h16 ;
            rom[14365] = 8'hec ;
            rom[14366] = 8'hd7 ;
            rom[14367] = 8'hf1 ;
            rom[14368] = 8'h0a ;
            rom[14369] = 8'he8 ;
            rom[14370] = 8'h17 ;
            rom[14371] = 8'hf4 ;
            rom[14372] = 8'hf4 ;
            rom[14373] = 8'h13 ;
            rom[14374] = 8'hb9 ;
            rom[14375] = 8'he0 ;
            rom[14376] = 8'h15 ;
            rom[14377] = 8'hff ;
            rom[14378] = 8'hff ;
            rom[14379] = 8'h0a ;
            rom[14380] = 8'hfb ;
            rom[14381] = 8'hf3 ;
            rom[14382] = 8'h0c ;
            rom[14383] = 8'h0a ;
            rom[14384] = 8'hec ;
            rom[14385] = 8'h1c ;
            rom[14386] = 8'hf5 ;
            rom[14387] = 8'he5 ;
            rom[14388] = 8'hf5 ;
            rom[14389] = 8'hef ;
            rom[14390] = 8'hee ;
            rom[14391] = 8'h06 ;
            rom[14392] = 8'hd7 ;
            rom[14393] = 8'h10 ;
            rom[14394] = 8'h09 ;
            rom[14395] = 8'hf1 ;
            rom[14396] = 8'he8 ;
            rom[14397] = 8'h0f ;
            rom[14398] = 8'hda ;
            rom[14399] = 8'he2 ;
            rom[14400] = 8'h0a ;
            rom[14401] = 8'hf5 ;
            rom[14402] = 8'h2b ;
            rom[14403] = 8'he3 ;
            rom[14404] = 8'heb ;
            rom[14405] = 8'hff ;
            rom[14406] = 8'h1f ;
            rom[14407] = 8'he1 ;
            rom[14408] = 8'he0 ;
            rom[14409] = 8'h22 ;
            rom[14410] = 8'h1e ;
            rom[14411] = 8'hf1 ;
            rom[14412] = 8'h03 ;
            rom[14413] = 8'h06 ;
            rom[14414] = 8'hec ;
            rom[14415] = 8'hda ;
            rom[14416] = 8'hf4 ;
            rom[14417] = 8'h10 ;
            rom[14418] = 8'h16 ;
            rom[14419] = 8'h08 ;
            rom[14420] = 8'h09 ;
            rom[14421] = 8'hea ;
            rom[14422] = 8'hf5 ;
            rom[14423] = 8'hfb ;
            rom[14424] = 8'he0 ;
            rom[14425] = 8'hbe ;
            rom[14426] = 8'hdb ;
            rom[14427] = 8'h08 ;
            rom[14428] = 8'hdd ;
            rom[14429] = 8'h06 ;
            rom[14430] = 8'h02 ;
            rom[14431] = 8'hf4 ;
            rom[14432] = 8'hf8 ;
            rom[14433] = 8'h05 ;
            rom[14434] = 8'hff ;
            rom[14435] = 8'h07 ;
            rom[14436] = 8'hdd ;
            rom[14437] = 8'hf3 ;
            rom[14438] = 8'h05 ;
            rom[14439] = 8'hfe ;
            rom[14440] = 8'hf6 ;
            rom[14441] = 8'h00 ;
            rom[14442] = 8'h07 ;
            rom[14443] = 8'h0d ;
            rom[14444] = 8'h15 ;
            rom[14445] = 8'h28 ;
            rom[14446] = 8'hf4 ;
            rom[14447] = 8'h10 ;
            rom[14448] = 8'hd4 ;
            rom[14449] = 8'he3 ;
            rom[14450] = 8'he5 ;
            rom[14451] = 8'hef ;
            rom[14452] = 8'hf3 ;
            rom[14453] = 8'h01 ;
            rom[14454] = 8'h18 ;
            rom[14455] = 8'h17 ;
            rom[14456] = 8'hfb ;
            rom[14457] = 8'hf0 ;
            rom[14458] = 8'hf1 ;
            rom[14459] = 8'h10 ;
            rom[14460] = 8'hfc ;
            rom[14461] = 8'h08 ;
            rom[14462] = 8'h13 ;
            rom[14463] = 8'h13 ;
            rom[14464] = 8'h02 ;
            rom[14465] = 8'h09 ;
            rom[14466] = 8'h0e ;
            rom[14467] = 8'h02 ;
            rom[14468] = 8'hed ;
            rom[14469] = 8'hd0 ;
            rom[14470] = 8'ha9 ;
            rom[14471] = 8'h1e ;
            rom[14472] = 8'h11 ;
            rom[14473] = 8'hc0 ;
            rom[14474] = 8'h03 ;
            rom[14475] = 8'hdf ;
            rom[14476] = 8'hf1 ;
            rom[14477] = 8'h02 ;
            rom[14478] = 8'h09 ;
            rom[14479] = 8'hd0 ;
            rom[14480] = 8'hf3 ;
            rom[14481] = 8'h07 ;
            rom[14482] = 8'hff ;
            rom[14483] = 8'h12 ;
            rom[14484] = 8'h0c ;
            rom[14485] = 8'h1f ;
            rom[14486] = 8'h27 ;
            rom[14487] = 8'hec ;
            rom[14488] = 8'he5 ;
            rom[14489] = 8'hff ;
            rom[14490] = 8'hdf ;
            rom[14491] = 8'hf1 ;
            rom[14492] = 8'he1 ;
            rom[14493] = 8'h0b ;
            rom[14494] = 8'hea ;
            rom[14495] = 8'h0f ;
            rom[14496] = 8'hf9 ;
            rom[14497] = 8'hea ;
            rom[14498] = 8'he8 ;
            rom[14499] = 8'he4 ;
            rom[14500] = 8'hfc ;
            rom[14501] = 8'h0b ;
            rom[14502] = 8'h07 ;
            rom[14503] = 8'hdc ;
            rom[14504] = 8'hf5 ;
            rom[14505] = 8'h06 ;
            rom[14506] = 8'hf9 ;
            rom[14507] = 8'h16 ;
            rom[14508] = 8'hfa ;
            rom[14509] = 8'hfa ;
            rom[14510] = 8'hf7 ;
            rom[14511] = 8'hfc ;
            rom[14512] = 8'h06 ;
            rom[14513] = 8'h18 ;
            rom[14514] = 8'h01 ;
            rom[14515] = 8'he4 ;
            rom[14516] = 8'h06 ;
            rom[14517] = 8'h1b ;
            rom[14518] = 8'hf0 ;
            rom[14519] = 8'hff ;
            rom[14520] = 8'hff ;
            rom[14521] = 8'h0b ;
            rom[14522] = 8'h17 ;
            rom[14523] = 8'hf8 ;
            rom[14524] = 8'h09 ;
            rom[14525] = 8'hd8 ;
            rom[14526] = 8'h1a ;
            rom[14527] = 8'he9 ;
            rom[14528] = 8'h13 ;
            rom[14529] = 8'h1f ;
            rom[14530] = 8'h09 ;
            rom[14531] = 8'hf0 ;
            rom[14532] = 8'hff ;
            rom[14533] = 8'he6 ;
            rom[14534] = 8'he7 ;
            rom[14535] = 8'h12 ;
            rom[14536] = 8'h02 ;
            rom[14537] = 8'heb ;
            rom[14538] = 8'h0b ;
            rom[14539] = 8'h0f ;
            rom[14540] = 8'hea ;
            rom[14541] = 8'h08 ;
            rom[14542] = 8'h22 ;
            rom[14543] = 8'hfc ;
            rom[14544] = 8'h0d ;
            rom[14545] = 8'hdb ;
            rom[14546] = 8'h08 ;
            rom[14547] = 8'hde ;
            rom[14548] = 8'hff ;
            rom[14549] = 8'h05 ;
            rom[14550] = 8'hd9 ;
            rom[14551] = 8'hcd ;
            rom[14552] = 8'h0b ;
            rom[14553] = 8'h12 ;
            rom[14554] = 8'h03 ;
            rom[14555] = 8'hf9 ;
            rom[14556] = 8'h1d ;
            rom[14557] = 8'hef ;
            rom[14558] = 8'h0f ;
            rom[14559] = 8'hf9 ;
            rom[14560] = 8'hf2 ;
            rom[14561] = 8'h13 ;
            rom[14562] = 8'h12 ;
            rom[14563] = 8'hfe ;
            rom[14564] = 8'hfc ;
            rom[14565] = 8'h08 ;
            rom[14566] = 8'he1 ;
            rom[14567] = 8'h0f ;
            rom[14568] = 8'hf0 ;
            rom[14569] = 8'h08 ;
            rom[14570] = 8'h0a ;
            rom[14571] = 8'h0b ;
            rom[14572] = 8'hf3 ;
            rom[14573] = 8'hd6 ;
            rom[14574] = 8'hf4 ;
            rom[14575] = 8'hd7 ;
            rom[14576] = 8'h1c ;
            rom[14577] = 8'h0f ;
            rom[14578] = 8'h04 ;
            rom[14579] = 8'hcd ;
            rom[14580] = 8'h10 ;
            rom[14581] = 8'hff ;
            rom[14582] = 8'h04 ;
            rom[14583] = 8'h20 ;
            rom[14584] = 8'h0d ;
            rom[14585] = 8'h04 ;
            rom[14586] = 8'h1c ;
            rom[14587] = 8'hfc ;
            rom[14588] = 8'hfd ;
            rom[14589] = 8'he6 ;
            rom[14590] = 8'hdf ;
            rom[14591] = 8'h03 ;
            rom[14592] = 8'h2d ;
            rom[14593] = 8'hf8 ;
            rom[14594] = 8'hfb ;
            rom[14595] = 8'h03 ;
            rom[14596] = 8'hfb ;
            rom[14597] = 8'h00 ;
            rom[14598] = 8'h29 ;
            rom[14599] = 8'h0c ;
            rom[14600] = 8'he9 ;
            rom[14601] = 8'h09 ;
            rom[14602] = 8'hfb ;
            rom[14603] = 8'hf2 ;
            rom[14604] = 8'he0 ;
            rom[14605] = 8'h10 ;
            rom[14606] = 8'h05 ;
            rom[14607] = 8'h08 ;
            rom[14608] = 8'hc0 ;
            rom[14609] = 8'hd0 ;
            rom[14610] = 8'h07 ;
            rom[14611] = 8'h0e ;
            rom[14612] = 8'hef ;
            rom[14613] = 8'he8 ;
            rom[14614] = 8'hd3 ;
            rom[14615] = 8'h15 ;
            rom[14616] = 8'h0e ;
            rom[14617] = 8'hed ;
            rom[14618] = 8'he7 ;
            rom[14619] = 8'hfd ;
            rom[14620] = 8'hfd ;
            rom[14621] = 8'h02 ;
            rom[14622] = 8'h02 ;
            rom[14623] = 8'h01 ;
            rom[14624] = 8'h0f ;
            rom[14625] = 8'hfd ;
            rom[14626] = 8'hf2 ;
            rom[14627] = 8'hca ;
            rom[14628] = 8'hfc ;
            rom[14629] = 8'hfe ;
            rom[14630] = 8'he9 ;
            rom[14631] = 8'hf9 ;
            rom[14632] = 8'hf4 ;
            rom[14633] = 8'h0f ;
            rom[14634] = 8'hf1 ;
            rom[14635] = 8'h0d ;
            rom[14636] = 8'hdf ;
            rom[14637] = 8'hf7 ;
            rom[14638] = 8'he7 ;
            rom[14639] = 8'hfc ;
            rom[14640] = 8'he7 ;
            rom[14641] = 8'h08 ;
            rom[14642] = 8'hf1 ;
            rom[14643] = 8'h10 ;
            rom[14644] = 8'h02 ;
            rom[14645] = 8'h03 ;
            rom[14646] = 8'he1 ;
            rom[14647] = 8'hdc ;
            rom[14648] = 8'h30 ;
            rom[14649] = 8'h0f ;
            rom[14650] = 8'h05 ;
            rom[14651] = 8'hf0 ;
            rom[14652] = 8'hff ;
            rom[14653] = 8'h0c ;
            rom[14654] = 8'hed ;
            rom[14655] = 8'h09 ;
            rom[14656] = 8'h0a ;
            rom[14657] = 8'hf4 ;
            rom[14658] = 8'hff ;
            rom[14659] = 8'h0c ;
            rom[14660] = 8'hf6 ;
            rom[14661] = 8'hfb ;
            rom[14662] = 8'hf7 ;
            rom[14663] = 8'h1a ;
            rom[14664] = 8'hef ;
            rom[14665] = 8'hfa ;
            rom[14666] = 8'h04 ;
            rom[14667] = 8'h05 ;
            rom[14668] = 8'hf7 ;
            rom[14669] = 8'h26 ;
            rom[14670] = 8'h00 ;
            rom[14671] = 8'hd4 ;
            rom[14672] = 8'hf8 ;
            rom[14673] = 8'h10 ;
            rom[14674] = 8'hff ;
            rom[14675] = 8'hdf ;
            rom[14676] = 8'h08 ;
            rom[14677] = 8'hda ;
            rom[14678] = 8'he7 ;
            rom[14679] = 8'h0f ;
            rom[14680] = 8'h15 ;
            rom[14681] = 8'hc5 ;
            rom[14682] = 8'h1c ;
            rom[14683] = 8'h08 ;
            rom[14684] = 8'h16 ;
            rom[14685] = 8'hf1 ;
            rom[14686] = 8'h09 ;
            rom[14687] = 8'h17 ;
            rom[14688] = 8'hff ;
            rom[14689] = 8'h02 ;
            rom[14690] = 8'hfb ;
            rom[14691] = 8'h05 ;
            rom[14692] = 8'h1b ;
            rom[14693] = 8'h03 ;
            rom[14694] = 8'hfb ;
            rom[14695] = 8'h23 ;
            rom[14696] = 8'hdc ;
            rom[14697] = 8'h07 ;
            rom[14698] = 8'he5 ;
            rom[14699] = 8'h13 ;
            rom[14700] = 8'h00 ;
            rom[14701] = 8'h04 ;
            rom[14702] = 8'h0e ;
            rom[14703] = 8'hea ;
            rom[14704] = 8'he5 ;
            rom[14705] = 8'h00 ;
            rom[14706] = 8'he6 ;
            rom[14707] = 8'h0f ;
            rom[14708] = 8'heb ;
            rom[14709] = 8'h0a ;
            rom[14710] = 8'hf1 ;
            rom[14711] = 8'hf4 ;
            rom[14712] = 8'hff ;
            rom[14713] = 8'h10 ;
            rom[14714] = 8'h0f ;
            rom[14715] = 8'h1d ;
            rom[14716] = 8'h20 ;
            rom[14717] = 8'hf1 ;
            rom[14718] = 8'h1a ;
            rom[14719] = 8'h08 ;
            rom[14720] = 8'hff ;
            rom[14721] = 8'hf7 ;
            rom[14722] = 8'h12 ;
            rom[14723] = 8'h07 ;
            rom[14724] = 8'hfd ;
            rom[14725] = 8'hc7 ;
            rom[14726] = 8'he1 ;
            rom[14727] = 8'h0d ;
            rom[14728] = 8'he8 ;
            rom[14729] = 8'he8 ;
            rom[14730] = 8'h13 ;
            rom[14731] = 8'h01 ;
            rom[14732] = 8'he0 ;
            rom[14733] = 8'h0a ;
            rom[14734] = 8'h1e ;
            rom[14735] = 8'h21 ;
            rom[14736] = 8'hf8 ;
            rom[14737] = 8'h21 ;
            rom[14738] = 8'h16 ;
            rom[14739] = 8'h0a ;
            rom[14740] = 8'h12 ;
            rom[14741] = 8'h03 ;
            rom[14742] = 8'h05 ;
            rom[14743] = 8'hfb ;
            rom[14744] = 8'hc8 ;
            rom[14745] = 8'h00 ;
            rom[14746] = 8'hf8 ;
            rom[14747] = 8'h0e ;
            rom[14748] = 8'hc2 ;
            rom[14749] = 8'h0e ;
            rom[14750] = 8'h01 ;
            rom[14751] = 8'h0e ;
            rom[14752] = 8'hd8 ;
            rom[14753] = 8'hf1 ;
            rom[14754] = 8'h03 ;
            rom[14755] = 8'hec ;
            rom[14756] = 8'h05 ;
            rom[14757] = 8'hf5 ;
            rom[14758] = 8'h04 ;
            rom[14759] = 8'hfa ;
            rom[14760] = 8'h12 ;
            rom[14761] = 8'hfc ;
            rom[14762] = 8'h0e ;
            rom[14763] = 8'hfb ;
            rom[14764] = 8'hfb ;
            rom[14765] = 8'hd4 ;
            rom[14766] = 8'he6 ;
            rom[14767] = 8'h06 ;
            rom[14768] = 8'h0a ;
            rom[14769] = 8'h06 ;
            rom[14770] = 8'hb0 ;
            rom[14771] = 8'hd3 ;
            rom[14772] = 8'h0d ;
            rom[14773] = 8'h07 ;
            rom[14774] = 8'hf4 ;
            rom[14775] = 8'hf9 ;
            rom[14776] = 8'hed ;
            rom[14777] = 8'h2d ;
            rom[14778] = 8'h02 ;
            rom[14779] = 8'h0a ;
            rom[14780] = 8'hdf ;
            rom[14781] = 8'hd0 ;
            rom[14782] = 8'h09 ;
            rom[14783] = 8'hf6 ;
            rom[14784] = 8'h2d ;
            rom[14785] = 8'h0c ;
            rom[14786] = 8'hee ;
            rom[14787] = 8'hfd ;
            rom[14788] = 8'hf3 ;
            rom[14789] = 8'h0f ;
            rom[14790] = 8'hfb ;
            rom[14791] = 8'h2a ;
            rom[14792] = 8'hf4 ;
            rom[14793] = 8'hf8 ;
            rom[14794] = 8'hf7 ;
            rom[14795] = 8'he7 ;
            rom[14796] = 8'hc4 ;
            rom[14797] = 8'he7 ;
            rom[14798] = 8'h10 ;
            rom[14799] = 8'hf3 ;
            rom[14800] = 8'h10 ;
            rom[14801] = 8'he1 ;
            rom[14802] = 8'h0a ;
            rom[14803] = 8'h02 ;
            rom[14804] = 8'hfd ;
            rom[14805] = 8'hf6 ;
            rom[14806] = 8'he9 ;
            rom[14807] = 8'h0b ;
            rom[14808] = 8'he5 ;
            rom[14809] = 8'hfd ;
            rom[14810] = 8'hf5 ;
            rom[14811] = 8'he4 ;
            rom[14812] = 8'hff ;
            rom[14813] = 8'hf2 ;
            rom[14814] = 8'h01 ;
            rom[14815] = 8'hf9 ;
            rom[14816] = 8'hd4 ;
            rom[14817] = 8'hdb ;
            rom[14818] = 8'h07 ;
            rom[14819] = 8'hfe ;
            rom[14820] = 8'h0f ;
            rom[14821] = 8'hfa ;
            rom[14822] = 8'h0d ;
            rom[14823] = 8'hf1 ;
            rom[14824] = 8'hf5 ;
            rom[14825] = 8'h14 ;
            rom[14826] = 8'he0 ;
            rom[14827] = 8'hff ;
            rom[14828] = 8'hc7 ;
            rom[14829] = 8'hf4 ;
            rom[14830] = 8'h01 ;
            rom[14831] = 8'hec ;
            rom[14832] = 8'h17 ;
            rom[14833] = 8'he8 ;
            rom[14834] = 8'hde ;
            rom[14835] = 8'hcf ;
            rom[14836] = 8'h0c ;
            rom[14837] = 8'h19 ;
            rom[14838] = 8'h03 ;
            rom[14839] = 8'h03 ;
            rom[14840] = 8'hff ;
            rom[14841] = 8'h10 ;
            rom[14842] = 8'h0e ;
            rom[14843] = 8'heb ;
            rom[14844] = 8'hee ;
            rom[14845] = 8'hcf ;
            rom[14846] = 8'h09 ;
            rom[14847] = 8'hfa ;
            rom[14848] = 8'h0a ;
            rom[14849] = 8'h13 ;
            rom[14850] = 8'h0f ;
            rom[14851] = 8'hed ;
            rom[14852] = 8'hdc ;
            rom[14853] = 8'h05 ;
            rom[14854] = 8'h1f ;
            rom[14855] = 8'he6 ;
            rom[14856] = 8'hde ;
            rom[14857] = 8'hfa ;
            rom[14858] = 8'h06 ;
            rom[14859] = 8'he1 ;
            rom[14860] = 8'hfc ;
            rom[14861] = 8'hfc ;
            rom[14862] = 8'hfa ;
            rom[14863] = 8'hf1 ;
            rom[14864] = 8'hcc ;
            rom[14865] = 8'h11 ;
            rom[14866] = 8'h0b ;
            rom[14867] = 8'hfc ;
            rom[14868] = 8'hce ;
            rom[14869] = 8'hce ;
            rom[14870] = 8'he8 ;
            rom[14871] = 8'h1d ;
            rom[14872] = 8'hfa ;
            rom[14873] = 8'h9c ;
            rom[14874] = 8'h09 ;
            rom[14875] = 8'hf9 ;
            rom[14876] = 8'h03 ;
            rom[14877] = 8'hfb ;
            rom[14878] = 8'h11 ;
            rom[14879] = 8'hf4 ;
            rom[14880] = 8'h18 ;
            rom[14881] = 8'hf0 ;
            rom[14882] = 8'hf4 ;
            rom[14883] = 8'hd6 ;
            rom[14884] = 8'hea ;
            rom[14885] = 8'h1b ;
            rom[14886] = 8'h05 ;
            rom[14887] = 8'h0b ;
            rom[14888] = 8'he6 ;
            rom[14889] = 8'hf7 ;
            rom[14890] = 8'hfc ;
            rom[14891] = 8'h08 ;
            rom[14892] = 8'h0d ;
            rom[14893] = 8'h04 ;
            rom[14894] = 8'hf1 ;
            rom[14895] = 8'he7 ;
            rom[14896] = 8'h20 ;
            rom[14897] = 8'hdb ;
            rom[14898] = 8'hec ;
            rom[14899] = 8'h03 ;
            rom[14900] = 8'hc7 ;
            rom[14901] = 8'h0c ;
            rom[14902] = 8'h12 ;
            rom[14903] = 8'hf4 ;
            rom[14904] = 8'h16 ;
            rom[14905] = 8'hfc ;
            rom[14906] = 8'h07 ;
            rom[14907] = 8'hfa ;
            rom[14908] = 8'h00 ;
            rom[14909] = 8'hf2 ;
            rom[14910] = 8'h0a ;
            rom[14911] = 8'hff ;
            rom[14912] = 8'h20 ;
            rom[14913] = 8'hef ;
            rom[14914] = 8'h18 ;
            rom[14915] = 8'hd7 ;
            rom[14916] = 8'hf9 ;
            rom[14917] = 8'h09 ;
            rom[14918] = 8'h10 ;
            rom[14919] = 8'hee ;
            rom[14920] = 8'hd4 ;
            rom[14921] = 8'hfd ;
            rom[14922] = 8'h0c ;
            rom[14923] = 8'he6 ;
            rom[14924] = 8'h0a ;
            rom[14925] = 8'hf7 ;
            rom[14926] = 8'hf3 ;
            rom[14927] = 8'he0 ;
            rom[14928] = 8'hdd ;
            rom[14929] = 8'h11 ;
            rom[14930] = 8'hf1 ;
            rom[14931] = 8'h0e ;
            rom[14932] = 8'h0b ;
            rom[14933] = 8'hcf ;
            rom[14934] = 8'hde ;
            rom[14935] = 8'h0f ;
            rom[14936] = 8'hf5 ;
            rom[14937] = 8'he9 ;
            rom[14938] = 8'heb ;
            rom[14939] = 8'h03 ;
            rom[14940] = 8'h1c ;
            rom[14941] = 8'hf6 ;
            rom[14942] = 8'h17 ;
            rom[14943] = 8'hf7 ;
            rom[14944] = 8'h04 ;
            rom[14945] = 8'hf0 ;
            rom[14946] = 8'hfc ;
            rom[14947] = 8'hd1 ;
            rom[14948] = 8'he2 ;
            rom[14949] = 8'h0f ;
            rom[14950] = 8'h0d ;
            rom[14951] = 8'hef ;
            rom[14952] = 8'hf5 ;
            rom[14953] = 8'hff ;
            rom[14954] = 8'hfe ;
            rom[14955] = 8'h14 ;
            rom[14956] = 8'h16 ;
            rom[14957] = 8'hfe ;
            rom[14958] = 8'h00 ;
            rom[14959] = 8'h11 ;
            rom[14960] = 8'hd7 ;
            rom[14961] = 8'hf7 ;
            rom[14962] = 8'hc7 ;
            rom[14963] = 8'hdd ;
            rom[14964] = 8'heb ;
            rom[14965] = 8'h0e ;
            rom[14966] = 8'h1f ;
            rom[14967] = 8'hf3 ;
            rom[14968] = 8'h06 ;
            rom[14969] = 8'h06 ;
            rom[14970] = 8'hfc ;
            rom[14971] = 8'hee ;
            rom[14972] = 8'hfe ;
            rom[14973] = 8'hfe ;
            rom[14974] = 8'h11 ;
            rom[14975] = 8'h06 ;
            rom[14976] = 8'he8 ;
            rom[14977] = 8'hf4 ;
            rom[14978] = 8'h0e ;
            rom[14979] = 8'h03 ;
            rom[14980] = 8'h18 ;
            rom[14981] = 8'hfd ;
            rom[14982] = 8'hed ;
            rom[14983] = 8'hfb ;
            rom[14984] = 8'h0d ;
            rom[14985] = 8'h16 ;
            rom[14986] = 8'hf4 ;
            rom[14987] = 8'h12 ;
            rom[14988] = 8'h13 ;
            rom[14989] = 8'h18 ;
            rom[14990] = 8'h17 ;
            rom[14991] = 8'hf8 ;
            rom[14992] = 8'hf5 ;
            rom[14993] = 8'h0b ;
            rom[14994] = 8'h0a ;
            rom[14995] = 8'h0c ;
            rom[14996] = 8'h15 ;
            rom[14997] = 8'heb ;
            rom[14998] = 8'hda ;
            rom[14999] = 8'hed ;
            rom[15000] = 8'h17 ;
            rom[15001] = 8'hf8 ;
            rom[15002] = 8'hf0 ;
            rom[15003] = 8'hdd ;
            rom[15004] = 8'h07 ;
            rom[15005] = 8'hfd ;
            rom[15006] = 8'h04 ;
            rom[15007] = 8'h0c ;
            rom[15008] = 8'hed ;
            rom[15009] = 8'hfd ;
            rom[15010] = 8'h13 ;
            rom[15011] = 8'hf0 ;
            rom[15012] = 8'h05 ;
            rom[15013] = 8'h0c ;
            rom[15014] = 8'h15 ;
            rom[15015] = 8'h03 ;
            rom[15016] = 8'hed ;
            rom[15017] = 8'h0b ;
            rom[15018] = 8'hea ;
            rom[15019] = 8'h0a ;
            rom[15020] = 8'h22 ;
            rom[15021] = 8'h0b ;
            rom[15022] = 8'h19 ;
            rom[15023] = 8'h12 ;
            rom[15024] = 8'hd3 ;
            rom[15025] = 8'h00 ;
            rom[15026] = 8'h16 ;
            rom[15027] = 8'hfc ;
            rom[15028] = 8'h0c ;
            rom[15029] = 8'h0b ;
            rom[15030] = 8'h03 ;
            rom[15031] = 8'hf3 ;
            rom[15032] = 8'h00 ;
            rom[15033] = 8'hf2 ;
            rom[15034] = 8'h06 ;
            rom[15035] = 8'h31 ;
            rom[15036] = 8'hfa ;
            rom[15037] = 8'h07 ;
            rom[15038] = 8'h05 ;
            rom[15039] = 8'he1 ;
            rom[15040] = 8'h13 ;
            rom[15041] = 8'h20 ;
            rom[15042] = 8'h11 ;
            rom[15043] = 8'h12 ;
            rom[15044] = 8'he3 ;
            rom[15045] = 8'hfb ;
            rom[15046] = 8'h09 ;
            rom[15047] = 8'hed ;
            rom[15048] = 8'heb ;
            rom[15049] = 8'hf5 ;
            rom[15050] = 8'hea ;
            rom[15051] = 8'h0b ;
            rom[15052] = 8'hfa ;
            rom[15053] = 8'h0b ;
            rom[15054] = 8'h09 ;
            rom[15055] = 8'hf6 ;
            rom[15056] = 8'hf5 ;
            rom[15057] = 8'hf9 ;
            rom[15058] = 8'h02 ;
            rom[15059] = 8'hd0 ;
            rom[15060] = 8'he7 ;
            rom[15061] = 8'hec ;
            rom[15062] = 8'h04 ;
            rom[15063] = 8'h04 ;
            rom[15064] = 8'h06 ;
            rom[15065] = 8'he8 ;
            rom[15066] = 8'hfa ;
            rom[15067] = 8'h02 ;
            rom[15068] = 8'h11 ;
            rom[15069] = 8'hf3 ;
            rom[15070] = 8'h0c ;
            rom[15071] = 8'h19 ;
            rom[15072] = 8'h1e ;
            rom[15073] = 8'hed ;
            rom[15074] = 8'he5 ;
            rom[15075] = 8'hf6 ;
            rom[15076] = 8'he0 ;
            rom[15077] = 8'h23 ;
            rom[15078] = 8'hf3 ;
            rom[15079] = 8'h0b ;
            rom[15080] = 8'hf0 ;
            rom[15081] = 8'hfc ;
            rom[15082] = 8'h15 ;
            rom[15083] = 8'h11 ;
            rom[15084] = 8'hfd ;
            rom[15085] = 8'h12 ;
            rom[15086] = 8'hf9 ;
            rom[15087] = 8'h1d ;
            rom[15088] = 8'hf5 ;
            rom[15089] = 8'h1a ;
            rom[15090] = 8'h0a ;
            rom[15091] = 8'h18 ;
            rom[15092] = 8'hec ;
            rom[15093] = 8'he1 ;
            rom[15094] = 8'hf7 ;
            rom[15095] = 8'h15 ;
            rom[15096] = 8'h16 ;
            rom[15097] = 8'hfe ;
            rom[15098] = 8'hfc ;
            rom[15099] = 8'hf4 ;
            rom[15100] = 8'hfe ;
            rom[15101] = 8'h15 ;
            rom[15102] = 8'hf2 ;
            rom[15103] = 8'h05 ;
            rom[15104] = 8'h0b ;
            rom[15105] = 8'hfb ;
            rom[15106] = 8'h12 ;
            rom[15107] = 8'he2 ;
            rom[15108] = 8'hfe ;
            rom[15109] = 8'hf0 ;
            rom[15110] = 8'hf1 ;
            rom[15111] = 8'hf4 ;
            rom[15112] = 8'hcf ;
            rom[15113] = 8'h08 ;
            rom[15114] = 8'h16 ;
            rom[15115] = 8'he2 ;
            rom[15116] = 8'hf7 ;
            rom[15117] = 8'hf4 ;
            rom[15118] = 8'he0 ;
            rom[15119] = 8'h0f ;
            rom[15120] = 8'hea ;
            rom[15121] = 8'h17 ;
            rom[15122] = 8'h06 ;
            rom[15123] = 8'h11 ;
            rom[15124] = 8'hfa ;
            rom[15125] = 8'h0b ;
            rom[15126] = 8'hfd ;
            rom[15127] = 8'h14 ;
            rom[15128] = 8'hcf ;
            rom[15129] = 8'hef ;
            rom[15130] = 8'had ;
            rom[15131] = 8'hfc ;
            rom[15132] = 8'hd6 ;
            rom[15133] = 8'h19 ;
            rom[15134] = 8'h0e ;
            rom[15135] = 8'hed ;
            rom[15136] = 8'h03 ;
            rom[15137] = 8'hf4 ;
            rom[15138] = 8'h11 ;
            rom[15139] = 8'h0d ;
            rom[15140] = 8'hfe ;
            rom[15141] = 8'hde ;
            rom[15142] = 8'hee ;
            rom[15143] = 8'hf6 ;
            rom[15144] = 8'h27 ;
            rom[15145] = 8'h03 ;
            rom[15146] = 8'hf6 ;
            rom[15147] = 8'h0a ;
            rom[15148] = 8'hf0 ;
            rom[15149] = 8'hef ;
            rom[15150] = 8'hee ;
            rom[15151] = 8'hdf ;
            rom[15152] = 8'hff ;
            rom[15153] = 8'h05 ;
            rom[15154] = 8'he0 ;
            rom[15155] = 8'hc4 ;
            rom[15156] = 8'h10 ;
            rom[15157] = 8'h0c ;
            rom[15158] = 8'h08 ;
            rom[15159] = 8'hfc ;
            rom[15160] = 8'hf7 ;
            rom[15161] = 8'hff ;
            rom[15162] = 8'he7 ;
            rom[15163] = 8'h17 ;
            rom[15164] = 8'hee ;
            rom[15165] = 8'hbb ;
            rom[15166] = 8'h2b ;
            rom[15167] = 8'hff ;
            rom[15168] = 8'h18 ;
            rom[15169] = 8'h01 ;
            rom[15170] = 8'h09 ;
            rom[15171] = 8'hf8 ;
            rom[15172] = 8'he1 ;
            rom[15173] = 8'hfa ;
            rom[15174] = 8'h1f ;
            rom[15175] = 8'hd8 ;
            rom[15176] = 8'he4 ;
            rom[15177] = 8'hff ;
            rom[15178] = 8'h12 ;
            rom[15179] = 8'h0d ;
            rom[15180] = 8'hb9 ;
            rom[15181] = 8'h0a ;
            rom[15182] = 8'he6 ;
            rom[15183] = 8'hea ;
            rom[15184] = 8'hf5 ;
            rom[15185] = 8'h00 ;
            rom[15186] = 8'hf1 ;
            rom[15187] = 8'hde ;
            rom[15188] = 8'he8 ;
            rom[15189] = 8'h08 ;
            rom[15190] = 8'h11 ;
            rom[15191] = 8'h1e ;
            rom[15192] = 8'h18 ;
            rom[15193] = 8'hf7 ;
            rom[15194] = 8'h10 ;
            rom[15195] = 8'he6 ;
            rom[15196] = 8'h03 ;
            rom[15197] = 8'h17 ;
            rom[15198] = 8'hfa ;
            rom[15199] = 8'h1a ;
            rom[15200] = 8'h1d ;
            rom[15201] = 8'h05 ;
            rom[15202] = 8'h11 ;
            rom[15203] = 8'h0f ;
            rom[15204] = 8'h07 ;
            rom[15205] = 8'h14 ;
            rom[15206] = 8'hdf ;
            rom[15207] = 8'h15 ;
            rom[15208] = 8'h12 ;
            rom[15209] = 8'h19 ;
            rom[15210] = 8'h1f ;
            rom[15211] = 8'hf9 ;
            rom[15212] = 8'hf9 ;
            rom[15213] = 8'h04 ;
            rom[15214] = 8'hfa ;
            rom[15215] = 8'hdf ;
            rom[15216] = 8'hff ;
            rom[15217] = 8'h15 ;
            rom[15218] = 8'h02 ;
            rom[15219] = 8'hf9 ;
            rom[15220] = 8'hb8 ;
            rom[15221] = 8'h02 ;
            rom[15222] = 8'hc5 ;
            rom[15223] = 8'h1e ;
            rom[15224] = 8'hf2 ;
            rom[15225] = 8'h19 ;
            rom[15226] = 8'hfb ;
            rom[15227] = 8'hed ;
            rom[15228] = 8'hf8 ;
            rom[15229] = 8'h12 ;
            rom[15230] = 8'he3 ;
            rom[15231] = 8'h14 ;
            rom[15232] = 8'h1e ;
            rom[15233] = 8'hf7 ;
            rom[15234] = 8'h00 ;
            rom[15235] = 8'hfd ;
            rom[15236] = 8'hee ;
            rom[15237] = 8'he7 ;
            rom[15238] = 8'hd8 ;
            rom[15239] = 8'heb ;
            rom[15240] = 8'hf2 ;
            rom[15241] = 8'hd0 ;
            rom[15242] = 8'h0e ;
            rom[15243] = 8'h16 ;
            rom[15244] = 8'hfe ;
            rom[15245] = 8'h1a ;
            rom[15246] = 8'h14 ;
            rom[15247] = 8'hf2 ;
            rom[15248] = 8'he2 ;
            rom[15249] = 8'h0e ;
            rom[15250] = 8'hec ;
            rom[15251] = 8'hf2 ;
            rom[15252] = 8'h11 ;
            rom[15253] = 8'h07 ;
            rom[15254] = 8'he7 ;
            rom[15255] = 8'hbb ;
            rom[15256] = 8'hef ;
            rom[15257] = 8'hfb ;
            rom[15258] = 8'hff ;
            rom[15259] = 8'he8 ;
            rom[15260] = 8'hfa ;
            rom[15261] = 8'hf8 ;
            rom[15262] = 8'hf6 ;
            rom[15263] = 8'hfc ;
            rom[15264] = 8'h1b ;
            rom[15265] = 8'hf5 ;
            rom[15266] = 8'h1f ;
            rom[15267] = 8'h01 ;
            rom[15268] = 8'he3 ;
            rom[15269] = 8'h15 ;
            rom[15270] = 8'hf1 ;
            rom[15271] = 8'hfb ;
            rom[15272] = 8'hf2 ;
            rom[15273] = 8'h05 ;
            rom[15274] = 8'h0a ;
            rom[15275] = 8'hee ;
            rom[15276] = 8'h19 ;
            rom[15277] = 8'h03 ;
            rom[15278] = 8'h0d ;
            rom[15279] = 8'h01 ;
            rom[15280] = 8'he3 ;
            rom[15281] = 8'h1d ;
            rom[15282] = 8'hd9 ;
            rom[15283] = 8'hf0 ;
            rom[15284] = 8'h07 ;
            rom[15285] = 8'h1c ;
            rom[15286] = 8'hfe ;
            rom[15287] = 8'hfb ;
            rom[15288] = 8'hf5 ;
            rom[15289] = 8'h02 ;
            rom[15290] = 8'h09 ;
            rom[15291] = 8'hf9 ;
            rom[15292] = 8'h06 ;
            rom[15293] = 8'hd7 ;
            rom[15294] = 8'hf6 ;
            rom[15295] = 8'hfa ;
            rom[15296] = 8'h07 ;
            rom[15297] = 8'he6 ;
            rom[15298] = 8'h18 ;
            rom[15299] = 8'hf5 ;
            rom[15300] = 8'hef ;
            rom[15301] = 8'h03 ;
            rom[15302] = 8'hf8 ;
            rom[15303] = 8'hff ;
            rom[15304] = 8'he0 ;
            rom[15305] = 8'h02 ;
            rom[15306] = 8'h09 ;
            rom[15307] = 8'h0a ;
            rom[15308] = 8'hf6 ;
            rom[15309] = 8'h0a ;
            rom[15310] = 8'hfd ;
            rom[15311] = 8'he2 ;
            rom[15312] = 8'hff ;
            rom[15313] = 8'hcd ;
            rom[15314] = 8'hec ;
            rom[15315] = 8'hee ;
            rom[15316] = 8'h0d ;
            rom[15317] = 8'h17 ;
            rom[15318] = 8'hf6 ;
            rom[15319] = 8'hfb ;
            rom[15320] = 8'he5 ;
            rom[15321] = 8'h02 ;
            rom[15322] = 8'hea ;
            rom[15323] = 8'h07 ;
            rom[15324] = 8'h0e ;
            rom[15325] = 8'h13 ;
            rom[15326] = 8'h20 ;
            rom[15327] = 8'hf3 ;
            rom[15328] = 8'h0f ;
            rom[15329] = 8'hf8 ;
            rom[15330] = 8'hff ;
            rom[15331] = 8'h03 ;
            rom[15332] = 8'he3 ;
            rom[15333] = 8'h21 ;
            rom[15334] = 8'hf4 ;
            rom[15335] = 8'hff ;
            rom[15336] = 8'h1f ;
            rom[15337] = 8'h02 ;
            rom[15338] = 8'hf8 ;
            rom[15339] = 8'h0a ;
            rom[15340] = 8'hee ;
            rom[15341] = 8'hf3 ;
            rom[15342] = 8'hfd ;
            rom[15343] = 8'hfc ;
            rom[15344] = 8'hce ;
            rom[15345] = 8'h0e ;
            rom[15346] = 8'hf5 ;
            rom[15347] = 8'hf0 ;
            rom[15348] = 8'h02 ;
            rom[15349] = 8'h2c ;
            rom[15350] = 8'h0e ;
            rom[15351] = 8'h16 ;
            rom[15352] = 8'h00 ;
            rom[15353] = 8'h14 ;
            rom[15354] = 8'h0c ;
            rom[15355] = 8'hdb ;
            rom[15356] = 8'hd4 ;
            rom[15357] = 8'h0c ;
            rom[15358] = 8'h23 ;
            rom[15359] = 8'h01 ;
            rom[15360] = 8'h05 ;
            rom[15361] = 8'h0c ;
            rom[15362] = 8'h17 ;
            rom[15363] = 8'hfd ;
            rom[15364] = 8'h09 ;
            rom[15365] = 8'hf4 ;
            rom[15366] = 8'hda ;
            rom[15367] = 8'h16 ;
            rom[15368] = 8'hfc ;
            rom[15369] = 8'h00 ;
            rom[15370] = 8'h0c ;
            rom[15371] = 8'hf9 ;
            rom[15372] = 8'h07 ;
            rom[15373] = 8'h14 ;
            rom[15374] = 8'hd7 ;
            rom[15375] = 8'h08 ;
            rom[15376] = 8'hfb ;
            rom[15377] = 8'he8 ;
            rom[15378] = 8'h0c ;
            rom[15379] = 8'hfe ;
            rom[15380] = 8'hf3 ;
            rom[15381] = 8'h05 ;
            rom[15382] = 8'hf1 ;
            rom[15383] = 8'he9 ;
            rom[15384] = 8'hee ;
            rom[15385] = 8'hfa ;
            rom[15386] = 8'hdf ;
            rom[15387] = 8'h11 ;
            rom[15388] = 8'hd5 ;
            rom[15389] = 8'h0a ;
            rom[15390] = 8'hfc ;
            rom[15391] = 8'h15 ;
            rom[15392] = 8'hdc ;
            rom[15393] = 8'h1c ;
            rom[15394] = 8'h05 ;
            rom[15395] = 8'h11 ;
            rom[15396] = 8'h01 ;
            rom[15397] = 8'hf0 ;
            rom[15398] = 8'h00 ;
            rom[15399] = 8'hd7 ;
            rom[15400] = 8'h15 ;
            rom[15401] = 8'hf6 ;
            rom[15402] = 8'h01 ;
            rom[15403] = 8'h06 ;
            rom[15404] = 8'h0c ;
            rom[15405] = 8'he6 ;
            rom[15406] = 8'hef ;
            rom[15407] = 8'h09 ;
            rom[15408] = 8'he8 ;
            rom[15409] = 8'hf8 ;
            rom[15410] = 8'hec ;
            rom[15411] = 8'hd1 ;
            rom[15412] = 8'h0b ;
            rom[15413] = 8'hfd ;
            rom[15414] = 8'h01 ;
            rom[15415] = 8'hf0 ;
            rom[15416] = 8'h0d ;
            rom[15417] = 8'h1d ;
            rom[15418] = 8'h04 ;
            rom[15419] = 8'hdf ;
            rom[15420] = 8'hde ;
            rom[15421] = 8'he0 ;
            rom[15422] = 8'h23 ;
            rom[15423] = 8'h07 ;
            rom[15424] = 8'hf9 ;
            rom[15425] = 8'h01 ;
            rom[15426] = 8'h19 ;
            rom[15427] = 8'he5 ;
            rom[15428] = 8'h0d ;
            rom[15429] = 8'h12 ;
            rom[15430] = 8'hfd ;
            rom[15431] = 8'h1d ;
            rom[15432] = 8'hf2 ;
            rom[15433] = 8'h15 ;
            rom[15434] = 8'hfd ;
            rom[15435] = 8'hc0 ;
            rom[15436] = 8'h03 ;
            rom[15437] = 8'he9 ;
            rom[15438] = 8'h15 ;
            rom[15439] = 8'h04 ;
            rom[15440] = 8'h0f ;
            rom[15441] = 8'hfe ;
            rom[15442] = 8'h21 ;
            rom[15443] = 8'hf1 ;
            rom[15444] = 8'he1 ;
            rom[15445] = 8'he9 ;
            rom[15446] = 8'h0d ;
            rom[15447] = 8'h01 ;
            rom[15448] = 8'hde ;
            rom[15449] = 8'hf2 ;
            rom[15450] = 8'h0d ;
            rom[15451] = 8'hd7 ;
            rom[15452] = 8'hfe ;
            rom[15453] = 8'h0c ;
            rom[15454] = 8'hc2 ;
            rom[15455] = 8'hfb ;
            rom[15456] = 8'h26 ;
            rom[15457] = 8'hde ;
            rom[15458] = 8'hf2 ;
            rom[15459] = 8'he0 ;
            rom[15460] = 8'h09 ;
            rom[15461] = 8'hfc ;
            rom[15462] = 8'h14 ;
            rom[15463] = 8'hf6 ;
            rom[15464] = 8'he4 ;
            rom[15465] = 8'h18 ;
            rom[15466] = 8'he6 ;
            rom[15467] = 8'h13 ;
            rom[15468] = 8'hdb ;
            rom[15469] = 8'h19 ;
            rom[15470] = 8'hf0 ;
            rom[15471] = 8'h11 ;
            rom[15472] = 8'h07 ;
            rom[15473] = 8'he9 ;
            rom[15474] = 8'h14 ;
            rom[15475] = 8'he0 ;
            rom[15476] = 8'h02 ;
            rom[15477] = 8'h0e ;
            rom[15478] = 8'h1a ;
            rom[15479] = 8'h15 ;
            rom[15480] = 8'hfc ;
            rom[15481] = 8'h08 ;
            rom[15482] = 8'h2a ;
            rom[15483] = 8'hee ;
            rom[15484] = 8'hf9 ;
            rom[15485] = 8'hec ;
            rom[15486] = 8'h01 ;
            rom[15487] = 8'he0 ;
            rom[15488] = 8'h09 ;
            rom[15489] = 8'h11 ;
            rom[15490] = 8'h14 ;
            rom[15491] = 8'hfc ;
            rom[15492] = 8'h15 ;
            rom[15493] = 8'h04 ;
            rom[15494] = 8'h02 ;
            rom[15495] = 8'hff ;
            rom[15496] = 8'hfd ;
            rom[15497] = 8'hff ;
            rom[15498] = 8'h20 ;
            rom[15499] = 8'h15 ;
            rom[15500] = 8'hc3 ;
            rom[15501] = 8'heb ;
            rom[15502] = 8'h0f ;
            rom[15503] = 8'h03 ;
            rom[15504] = 8'h08 ;
            rom[15505] = 8'hf2 ;
            rom[15506] = 8'h28 ;
            rom[15507] = 8'h0e ;
            rom[15508] = 8'he8 ;
            rom[15509] = 8'h03 ;
            rom[15510] = 8'hfd ;
            rom[15511] = 8'h0e ;
            rom[15512] = 8'hda ;
            rom[15513] = 8'hfe ;
            rom[15514] = 8'hcf ;
            rom[15515] = 8'h01 ;
            rom[15516] = 8'hb6 ;
            rom[15517] = 8'h0b ;
            rom[15518] = 8'h06 ;
            rom[15519] = 8'h04 ;
            rom[15520] = 8'hf5 ;
            rom[15521] = 8'h02 ;
            rom[15522] = 8'h06 ;
            rom[15523] = 8'hf0 ;
            rom[15524] = 8'h18 ;
            rom[15525] = 8'hfd ;
            rom[15526] = 8'hfa ;
            rom[15527] = 8'h01 ;
            rom[15528] = 8'h2d ;
            rom[15529] = 8'h03 ;
            rom[15530] = 8'h0a ;
            rom[15531] = 8'hfc ;
            rom[15532] = 8'hc7 ;
            rom[15533] = 8'hbb ;
            rom[15534] = 8'h04 ;
            rom[15535] = 8'hf6 ;
            rom[15536] = 8'h00 ;
            rom[15537] = 8'h03 ;
            rom[15538] = 8'he3 ;
            rom[15539] = 8'hec ;
            rom[15540] = 8'hef ;
            rom[15541] = 8'h0f ;
            rom[15542] = 8'hfa ;
            rom[15543] = 8'hed ;
            rom[15544] = 8'h00 ;
            rom[15545] = 8'h07 ;
            rom[15546] = 8'he5 ;
            rom[15547] = 8'h18 ;
            rom[15548] = 8'hd6 ;
            rom[15549] = 8'hd5 ;
            rom[15550] = 8'h0f ;
            rom[15551] = 8'hf8 ;
            rom[15552] = 8'h06 ;
            rom[15553] = 8'h14 ;
            rom[15554] = 8'hee ;
            rom[15555] = 8'h1c ;
            rom[15556] = 8'hc5 ;
            rom[15557] = 8'hc8 ;
            rom[15558] = 8'h05 ;
            rom[15559] = 8'h02 ;
            rom[15560] = 8'hf3 ;
            rom[15561] = 8'h0d ;
            rom[15562] = 8'he9 ;
            rom[15563] = 8'hff ;
            rom[15564] = 8'hfc ;
            rom[15565] = 8'h0d ;
            rom[15566] = 8'hee ;
            rom[15567] = 8'hf5 ;
            rom[15568] = 8'hc4 ;
            rom[15569] = 8'he1 ;
            rom[15570] = 8'h0e ;
            rom[15571] = 8'heb ;
            rom[15572] = 8'h19 ;
            rom[15573] = 8'hff ;
            rom[15574] = 8'hf6 ;
            rom[15575] = 8'hea ;
            rom[15576] = 8'h1e ;
            rom[15577] = 8'hd5 ;
            rom[15578] = 8'hff ;
            rom[15579] = 8'hea ;
            rom[15580] = 8'h13 ;
            rom[15581] = 8'hff ;
            rom[15582] = 8'hfc ;
            rom[15583] = 8'hed ;
            rom[15584] = 8'h1a ;
            rom[15585] = 8'he3 ;
            rom[15586] = 8'h1c ;
            rom[15587] = 8'hce ;
            rom[15588] = 8'hf3 ;
            rom[15589] = 8'h06 ;
            rom[15590] = 8'h00 ;
            rom[15591] = 8'h01 ;
            rom[15592] = 8'h06 ;
            rom[15593] = 8'hde ;
            rom[15594] = 8'hc5 ;
            rom[15595] = 8'h3a ;
            rom[15596] = 8'hf1 ;
            rom[15597] = 8'h0b ;
            rom[15598] = 8'hcd ;
            rom[15599] = 8'hff ;
            rom[15600] = 8'h1e ;
            rom[15601] = 8'hd8 ;
            rom[15602] = 8'h0e ;
            rom[15603] = 8'h0a ;
            rom[15604] = 8'he5 ;
            rom[15605] = 8'h00 ;
            rom[15606] = 8'hc6 ;
            rom[15607] = 8'h09 ;
            rom[15608] = 8'h0b ;
            rom[15609] = 8'h0d ;
            rom[15610] = 8'hf8 ;
            rom[15611] = 8'h14 ;
            rom[15612] = 8'h15 ;
            rom[15613] = 8'hfd ;
            rom[15614] = 8'h1a ;
            rom[15615] = 8'h06 ;
            rom[15616] = 8'h26 ;
            rom[15617] = 8'h05 ;
            rom[15618] = 8'h0b ;
            rom[15619] = 8'hf7 ;
            rom[15620] = 8'h02 ;
            rom[15621] = 8'h0e ;
            rom[15622] = 8'h19 ;
            rom[15623] = 8'h00 ;
            rom[15624] = 8'h07 ;
            rom[15625] = 8'hff ;
            rom[15626] = 8'h16 ;
            rom[15627] = 8'hfe ;
            rom[15628] = 8'h0e ;
            rom[15629] = 8'h22 ;
            rom[15630] = 8'he0 ;
            rom[15631] = 8'hf5 ;
            rom[15632] = 8'hfc ;
            rom[15633] = 8'hff ;
            rom[15634] = 8'h00 ;
            rom[15635] = 8'h0c ;
            rom[15636] = 8'hfe ;
            rom[15637] = 8'hd3 ;
            rom[15638] = 8'hf3 ;
            rom[15639] = 8'h0a ;
            rom[15640] = 8'he1 ;
            rom[15641] = 8'hd3 ;
            rom[15642] = 8'he5 ;
            rom[15643] = 8'h10 ;
            rom[15644] = 8'hf4 ;
            rom[15645] = 8'heb ;
            rom[15646] = 8'hee ;
            rom[15647] = 8'h05 ;
            rom[15648] = 8'hee ;
            rom[15649] = 8'h12 ;
            rom[15650] = 8'h0d ;
            rom[15651] = 8'hfd ;
            rom[15652] = 8'h03 ;
            rom[15653] = 8'hfe ;
            rom[15654] = 8'hd4 ;
            rom[15655] = 8'hde ;
            rom[15656] = 8'h0b ;
            rom[15657] = 8'h0a ;
            rom[15658] = 8'h00 ;
            rom[15659] = 8'h08 ;
            rom[15660] = 8'h01 ;
            rom[15661] = 8'h05 ;
            rom[15662] = 8'hf4 ;
            rom[15663] = 8'h02 ;
            rom[15664] = 8'he9 ;
            rom[15665] = 8'h0f ;
            rom[15666] = 8'hd2 ;
            rom[15667] = 8'hf9 ;
            rom[15668] = 8'hf1 ;
            rom[15669] = 8'hf7 ;
            rom[15670] = 8'h17 ;
            rom[15671] = 8'he2 ;
            rom[15672] = 8'h0f ;
            rom[15673] = 8'h08 ;
            rom[15674] = 8'he7 ;
            rom[15675] = 8'hfd ;
            rom[15676] = 8'hfc ;
            rom[15677] = 8'hf6 ;
            rom[15678] = 8'h04 ;
            rom[15679] = 8'h0b ;
            rom[15680] = 8'h08 ;
            rom[15681] = 8'h11 ;
            rom[15682] = 8'h12 ;
            rom[15683] = 8'h0f ;
            rom[15684] = 8'hfe ;
            rom[15685] = 8'hdb ;
            rom[15686] = 8'hbf ;
            rom[15687] = 8'h07 ;
            rom[15688] = 8'hff ;
            rom[15689] = 8'h03 ;
            rom[15690] = 8'hf7 ;
            rom[15691] = 8'h0b ;
            rom[15692] = 8'h0f ;
            rom[15693] = 8'h10 ;
            rom[15694] = 8'h0b ;
            rom[15695] = 8'hdc ;
            rom[15696] = 8'hf4 ;
            rom[15697] = 8'hfb ;
            rom[15698] = 8'h22 ;
            rom[15699] = 8'h00 ;
            rom[15700] = 8'h06 ;
            rom[15701] = 8'he9 ;
            rom[15702] = 8'hef ;
            rom[15703] = 8'h0a ;
            rom[15704] = 8'hfe ;
            rom[15705] = 8'h04 ;
            rom[15706] = 8'he4 ;
            rom[15707] = 8'hfe ;
            rom[15708] = 8'h03 ;
            rom[15709] = 8'hef ;
            rom[15710] = 8'hee ;
            rom[15711] = 8'h16 ;
            rom[15712] = 8'h19 ;
            rom[15713] = 8'h02 ;
            rom[15714] = 8'hf8 ;
            rom[15715] = 8'h13 ;
            rom[15716] = 8'h0a ;
            rom[15717] = 8'hf6 ;
            rom[15718] = 8'hf9 ;
            rom[15719] = 8'hdb ;
            rom[15720] = 8'heb ;
            rom[15721] = 8'hd4 ;
            rom[15722] = 8'h00 ;
            rom[15723] = 8'h1c ;
            rom[15724] = 8'h0d ;
            rom[15725] = 8'hed ;
            rom[15726] = 8'he7 ;
            rom[15727] = 8'h04 ;
            rom[15728] = 8'hfd ;
            rom[15729] = 8'h04 ;
            rom[15730] = 8'h04 ;
            rom[15731] = 8'h00 ;
            rom[15732] = 8'hfd ;
            rom[15733] = 8'hff ;
            rom[15734] = 8'hfb ;
            rom[15735] = 8'h04 ;
            rom[15736] = 8'heb ;
            rom[15737] = 8'hf7 ;
            rom[15738] = 8'h1b ;
            rom[15739] = 8'hf3 ;
            rom[15740] = 8'h23 ;
            rom[15741] = 8'h0d ;
            rom[15742] = 8'h28 ;
            rom[15743] = 8'hf5 ;
            rom[15744] = 8'h17 ;
            rom[15745] = 8'hf1 ;
            rom[15746] = 8'heb ;
            rom[15747] = 8'h12 ;
            rom[15748] = 8'hf3 ;
            rom[15749] = 8'h0b ;
            rom[15750] = 8'h07 ;
            rom[15751] = 8'h01 ;
            rom[15752] = 8'hf9 ;
            rom[15753] = 8'h0a ;
            rom[15754] = 8'h03 ;
            rom[15755] = 8'h12 ;
            rom[15756] = 8'heb ;
            rom[15757] = 8'hf0 ;
            rom[15758] = 8'hf9 ;
            rom[15759] = 8'hcd ;
            rom[15760] = 8'hf6 ;
            rom[15761] = 8'h05 ;
            rom[15762] = 8'hfe ;
            rom[15763] = 8'he0 ;
            rom[15764] = 8'hf3 ;
            rom[15765] = 8'hfd ;
            rom[15766] = 8'he5 ;
            rom[15767] = 8'h01 ;
            rom[15768] = 8'h15 ;
            rom[15769] = 8'hd6 ;
            rom[15770] = 8'hf8 ;
            rom[15771] = 8'hf6 ;
            rom[15772] = 8'hf2 ;
            rom[15773] = 8'hf1 ;
            rom[15774] = 8'hf9 ;
            rom[15775] = 8'h10 ;
            rom[15776] = 8'h1d ;
            rom[15777] = 8'hf6 ;
            rom[15778] = 8'hf3 ;
            rom[15779] = 8'hf6 ;
            rom[15780] = 8'hf9 ;
            rom[15781] = 8'hfa ;
            rom[15782] = 8'h0a ;
            rom[15783] = 8'h1b ;
            rom[15784] = 8'hd5 ;
            rom[15785] = 8'hfa ;
            rom[15786] = 8'hf6 ;
            rom[15787] = 8'h02 ;
            rom[15788] = 8'he6 ;
            rom[15789] = 8'h00 ;
            rom[15790] = 8'h19 ;
            rom[15791] = 8'hbf ;
            rom[15792] = 8'hef ;
            rom[15793] = 8'hfe ;
            rom[15794] = 8'hcd ;
            rom[15795] = 8'h00 ;
            rom[15796] = 8'hcb ;
            rom[15797] = 8'hf4 ;
            rom[15798] = 8'h05 ;
            rom[15799] = 8'h01 ;
            rom[15800] = 8'hf8 ;
            rom[15801] = 8'hf3 ;
            rom[15802] = 8'h19 ;
            rom[15803] = 8'h10 ;
            rom[15804] = 8'h24 ;
            rom[15805] = 8'hec ;
            rom[15806] = 8'h10 ;
            rom[15807] = 8'h1a ;
            rom[15808] = 8'h03 ;
            rom[15809] = 8'h0d ;
            rom[15810] = 8'h2a ;
            rom[15811] = 8'hee ;
            rom[15812] = 8'h02 ;
            rom[15813] = 8'h06 ;
            rom[15814] = 8'hf3 ;
            rom[15815] = 8'h19 ;
            rom[15816] = 8'h01 ;
            rom[15817] = 8'h00 ;
            rom[15818] = 8'h04 ;
            rom[15819] = 8'h28 ;
            rom[15820] = 8'he5 ;
            rom[15821] = 8'h00 ;
            rom[15822] = 8'h07 ;
            rom[15823] = 8'hd7 ;
            rom[15824] = 8'hd6 ;
            rom[15825] = 8'h02 ;
            rom[15826] = 8'h12 ;
            rom[15827] = 8'h0c ;
            rom[15828] = 8'hf2 ;
            rom[15829] = 8'hed ;
            rom[15830] = 8'h0b ;
            rom[15831] = 8'hf9 ;
            rom[15832] = 8'hf8 ;
            rom[15833] = 8'h0b ;
            rom[15834] = 8'hef ;
            rom[15835] = 8'he9 ;
            rom[15836] = 8'he5 ;
            rom[15837] = 8'he3 ;
            rom[15838] = 8'hcb ;
            rom[15839] = 8'hff ;
            rom[15840] = 8'hf0 ;
            rom[15841] = 8'hf7 ;
            rom[15842] = 8'h0d ;
            rom[15843] = 8'hf4 ;
            rom[15844] = 8'h19 ;
            rom[15845] = 8'hec ;
            rom[15846] = 8'h0e ;
            rom[15847] = 8'he6 ;
            rom[15848] = 8'hfb ;
            rom[15849] = 8'hfd ;
            rom[15850] = 8'h14 ;
            rom[15851] = 8'h10 ;
            rom[15852] = 8'h05 ;
            rom[15853] = 8'h01 ;
            rom[15854] = 8'h0a ;
            rom[15855] = 8'h23 ;
            rom[15856] = 8'he9 ;
            rom[15857] = 8'h0f ;
            rom[15858] = 8'h09 ;
            rom[15859] = 8'h12 ;
            rom[15860] = 8'hd6 ;
            rom[15861] = 8'h08 ;
            rom[15862] = 8'hec ;
            rom[15863] = 8'hfd ;
            rom[15864] = 8'hfb ;
            rom[15865] = 8'hf1 ;
            rom[15866] = 8'h06 ;
            rom[15867] = 8'h09 ;
            rom[15868] = 8'h27 ;
            rom[15869] = 8'h0c ;
            rom[15870] = 8'h05 ;
            rom[15871] = 8'h0c ;
            rom[15872] = 8'h2c ;
            rom[15873] = 8'hd1 ;
            rom[15874] = 8'h09 ;
            rom[15875] = 8'hf8 ;
            rom[15876] = 8'h02 ;
            rom[15877] = 8'h0e ;
            rom[15878] = 8'h10 ;
            rom[15879] = 8'h12 ;
            rom[15880] = 8'hdc ;
            rom[15881] = 8'h0b ;
            rom[15882] = 8'h10 ;
            rom[15883] = 8'hfa ;
            rom[15884] = 8'hf1 ;
            rom[15885] = 8'hfe ;
            rom[15886] = 8'he5 ;
            rom[15887] = 8'he9 ;
            rom[15888] = 8'hf7 ;
            rom[15889] = 8'h03 ;
            rom[15890] = 8'h18 ;
            rom[15891] = 8'h10 ;
            rom[15892] = 8'he5 ;
            rom[15893] = 8'h06 ;
            rom[15894] = 8'hf6 ;
            rom[15895] = 8'h06 ;
            rom[15896] = 8'hfd ;
            rom[15897] = 8'hdd ;
            rom[15898] = 8'he2 ;
            rom[15899] = 8'hd6 ;
            rom[15900] = 8'hf0 ;
            rom[15901] = 8'hed ;
            rom[15902] = 8'h09 ;
            rom[15903] = 8'hff ;
            rom[15904] = 8'hfb ;
            rom[15905] = 8'he2 ;
            rom[15906] = 8'hed ;
            rom[15907] = 8'hf8 ;
            rom[15908] = 8'hf7 ;
            rom[15909] = 8'hf0 ;
            rom[15910] = 8'h00 ;
            rom[15911] = 8'hf4 ;
            rom[15912] = 8'h00 ;
            rom[15913] = 8'h10 ;
            rom[15914] = 8'h0f ;
            rom[15915] = 8'h0f ;
            rom[15916] = 8'hfa ;
            rom[15917] = 8'h1b ;
            rom[15918] = 8'hf7 ;
            rom[15919] = 8'h0a ;
            rom[15920] = 8'hfb ;
            rom[15921] = 8'hef ;
            rom[15922] = 8'hf3 ;
            rom[15923] = 8'hd2 ;
            rom[15924] = 8'hef ;
            rom[15925] = 8'h1b ;
            rom[15926] = 8'h17 ;
            rom[15927] = 8'hf0 ;
            rom[15928] = 8'h07 ;
            rom[15929] = 8'hed ;
            rom[15930] = 8'h00 ;
            rom[15931] = 8'h09 ;
            rom[15932] = 8'h15 ;
            rom[15933] = 8'hef ;
            rom[15934] = 8'h11 ;
            rom[15935] = 8'h23 ;
            rom[15936] = 8'hf2 ;
            rom[15937] = 8'h13 ;
            rom[15938] = 8'h01 ;
            rom[15939] = 8'h12 ;
            rom[15940] = 8'hb1 ;
            rom[15941] = 8'hf8 ;
            rom[15942] = 8'hf6 ;
            rom[15943] = 8'hf9 ;
            rom[15944] = 8'hc6 ;
            rom[15945] = 8'h15 ;
            rom[15946] = 8'hf9 ;
            rom[15947] = 8'hed ;
            rom[15948] = 8'hf0 ;
            rom[15949] = 8'h0a ;
            rom[15950] = 8'h06 ;
            rom[15951] = 8'h02 ;
            rom[15952] = 8'ha7 ;
            rom[15953] = 8'hf8 ;
            rom[15954] = 8'h1a ;
            rom[15955] = 8'hff ;
            rom[15956] = 8'he5 ;
            rom[15957] = 8'hfa ;
            rom[15958] = 8'he6 ;
            rom[15959] = 8'he5 ;
            rom[15960] = 8'h16 ;
            rom[15961] = 8'hba ;
            rom[15962] = 8'h03 ;
            rom[15963] = 8'hf8 ;
            rom[15964] = 8'hf3 ;
            rom[15965] = 8'he4 ;
            rom[15966] = 8'h02 ;
            rom[15967] = 8'hf6 ;
            rom[15968] = 8'h2b ;
            rom[15969] = 8'hee ;
            rom[15970] = 8'h1a ;
            rom[15971] = 8'hdf ;
            rom[15972] = 8'he1 ;
            rom[15973] = 8'hf7 ;
            rom[15974] = 8'h04 ;
            rom[15975] = 8'hfc ;
            rom[15976] = 8'hf0 ;
            rom[15977] = 8'hec ;
            rom[15978] = 8'he5 ;
            rom[15979] = 8'h27 ;
            rom[15980] = 8'hf0 ;
            rom[15981] = 8'hff ;
            rom[15982] = 8'hd8 ;
            rom[15983] = 8'h02 ;
            rom[15984] = 8'h14 ;
            rom[15985] = 8'h05 ;
            rom[15986] = 8'he9 ;
            rom[15987] = 8'h06 ;
            rom[15988] = 8'hc8 ;
            rom[15989] = 8'hf0 ;
            rom[15990] = 8'hda ;
            rom[15991] = 8'h02 ;
            rom[15992] = 8'h0b ;
            rom[15993] = 8'hf5 ;
            rom[15994] = 8'h02 ;
            rom[15995] = 8'h0c ;
            rom[15996] = 8'h06 ;
            rom[15997] = 8'h0e ;
            rom[15998] = 8'h1b ;
            rom[15999] = 8'hf9 ;
            rom[16000] = 8'hf2 ;
            rom[16001] = 8'h15 ;
            rom[16002] = 8'hf9 ;
            rom[16003] = 8'h1a ;
            rom[16004] = 8'hae ;
            rom[16005] = 8'hde ;
            rom[16006] = 8'hfb ;
            rom[16007] = 8'h02 ;
            rom[16008] = 8'hd0 ;
            rom[16009] = 8'hf7 ;
            rom[16010] = 8'hf7 ;
            rom[16011] = 8'hf0 ;
            rom[16012] = 8'hfb ;
            rom[16013] = 8'h11 ;
            rom[16014] = 8'h00 ;
            rom[16015] = 8'hf1 ;
            rom[16016] = 8'hc7 ;
            rom[16017] = 8'h09 ;
            rom[16018] = 8'h19 ;
            rom[16019] = 8'hd9 ;
            rom[16020] = 8'hce ;
            rom[16021] = 8'hcc ;
            rom[16022] = 8'hff ;
            rom[16023] = 8'h08 ;
            rom[16024] = 8'h0c ;
            rom[16025] = 8'ha8 ;
            rom[16026] = 8'h09 ;
            rom[16027] = 8'hf0 ;
            rom[16028] = 8'h0b ;
            rom[16029] = 8'hfe ;
            rom[16030] = 8'h0d ;
            rom[16031] = 8'he9 ;
            rom[16032] = 8'h13 ;
            rom[16033] = 8'hc6 ;
            rom[16034] = 8'h05 ;
            rom[16035] = 8'hd0 ;
            rom[16036] = 8'hea ;
            rom[16037] = 8'h09 ;
            rom[16038] = 8'h16 ;
            rom[16039] = 8'h0e ;
            rom[16040] = 8'he6 ;
            rom[16041] = 8'h05 ;
            rom[16042] = 8'hfd ;
            rom[16043] = 8'h16 ;
            rom[16044] = 8'h03 ;
            rom[16045] = 8'h15 ;
            rom[16046] = 8'hf3 ;
            rom[16047] = 8'hdc ;
            rom[16048] = 8'h2f ;
            rom[16049] = 8'hfa ;
            rom[16050] = 8'hf2 ;
            rom[16051] = 8'h0f ;
            rom[16052] = 8'hcb ;
            rom[16053] = 8'hfb ;
            rom[16054] = 8'hfc ;
            rom[16055] = 8'hed ;
            rom[16056] = 8'h16 ;
            rom[16057] = 8'hf4 ;
            rom[16058] = 8'h1b ;
            rom[16059] = 8'h02 ;
            rom[16060] = 8'h19 ;
            rom[16061] = 8'hfd ;
            rom[16062] = 8'h04 ;
            rom[16063] = 8'hee ;
            rom[16064] = 8'h09 ;
            rom[16065] = 8'h05 ;
            rom[16066] = 8'h1a ;
            rom[16067] = 8'h0d ;
            rom[16068] = 8'hef ;
            rom[16069] = 8'hd9 ;
            rom[16070] = 8'he1 ;
            rom[16071] = 8'h08 ;
            rom[16072] = 8'hf4 ;
            rom[16073] = 8'h09 ;
            rom[16074] = 8'h04 ;
            rom[16075] = 8'h26 ;
            rom[16076] = 8'h0a ;
            rom[16077] = 8'hff ;
            rom[16078] = 8'hf5 ;
            rom[16079] = 8'hf7 ;
            rom[16080] = 8'hbe ;
            rom[16081] = 8'hf0 ;
            rom[16082] = 8'h1b ;
            rom[16083] = 8'hf2 ;
            rom[16084] = 8'hee ;
            rom[16085] = 8'hf5 ;
            rom[16086] = 8'h0d ;
            rom[16087] = 8'hf1 ;
            rom[16088] = 8'h0e ;
            rom[16089] = 8'he1 ;
            rom[16090] = 8'h1b ;
            rom[16091] = 8'hd3 ;
            rom[16092] = 8'hfc ;
            rom[16093] = 8'he1 ;
            rom[16094] = 8'he6 ;
            rom[16095] = 8'h13 ;
            rom[16096] = 8'h0a ;
            rom[16097] = 8'hfe ;
            rom[16098] = 8'hfa ;
            rom[16099] = 8'hc6 ;
            rom[16100] = 8'h1b ;
            rom[16101] = 8'h07 ;
            rom[16102] = 8'h04 ;
            rom[16103] = 8'h04 ;
            rom[16104] = 8'hfb ;
            rom[16105] = 8'he4 ;
            rom[16106] = 8'h05 ;
            rom[16107] = 8'h25 ;
            rom[16108] = 8'h09 ;
            rom[16109] = 8'h00 ;
            rom[16110] = 8'h19 ;
            rom[16111] = 8'hfc ;
            rom[16112] = 8'h0d ;
            rom[16113] = 8'h09 ;
            rom[16114] = 8'hf0 ;
            rom[16115] = 8'h17 ;
            rom[16116] = 8'he9 ;
            rom[16117] = 8'hfa ;
            rom[16118] = 8'hd3 ;
            rom[16119] = 8'h0a ;
            rom[16120] = 8'h0c ;
            rom[16121] = 8'h0e ;
            rom[16122] = 8'h19 ;
            rom[16123] = 8'h03 ;
            rom[16124] = 8'h1b ;
            rom[16125] = 8'h14 ;
            rom[16126] = 8'h04 ;
            rom[16127] = 8'h0a ;
            rom[16128] = 8'hf8 ;
            rom[16129] = 8'h07 ;
            rom[16130] = 8'h29 ;
            rom[16131] = 8'h13 ;
            rom[16132] = 8'hf4 ;
            rom[16133] = 8'h01 ;
            rom[16134] = 8'hdd ;
            rom[16135] = 8'hf6 ;
            rom[16136] = 8'hef ;
            rom[16137] = 8'h0b ;
            rom[16138] = 8'h04 ;
            rom[16139] = 8'hfe ;
            rom[16140] = 8'h05 ;
            rom[16141] = 8'h0d ;
            rom[16142] = 8'hef ;
            rom[16143] = 8'heb ;
            rom[16144] = 8'h02 ;
            rom[16145] = 8'h17 ;
            rom[16146] = 8'h03 ;
            rom[16147] = 8'h05 ;
            rom[16148] = 8'h1e ;
            rom[16149] = 8'hf5 ;
            rom[16150] = 8'hbc ;
            rom[16151] = 8'hf3 ;
            rom[16152] = 8'hed ;
            rom[16153] = 8'hed ;
            rom[16154] = 8'h14 ;
            rom[16155] = 8'h04 ;
            rom[16156] = 8'he4 ;
            rom[16157] = 8'he9 ;
            rom[16158] = 8'he9 ;
            rom[16159] = 8'h13 ;
            rom[16160] = 8'hf1 ;
            rom[16161] = 8'h0a ;
            rom[16162] = 8'h15 ;
            rom[16163] = 8'h20 ;
            rom[16164] = 8'h08 ;
            rom[16165] = 8'hf3 ;
            rom[16166] = 8'hed ;
            rom[16167] = 8'hfd ;
            rom[16168] = 8'hf6 ;
            rom[16169] = 8'hf8 ;
            rom[16170] = 8'hfc ;
            rom[16171] = 8'hdb ;
            rom[16172] = 8'h04 ;
            rom[16173] = 8'he3 ;
            rom[16174] = 8'h0e ;
            rom[16175] = 8'h1a ;
            rom[16176] = 8'hea ;
            rom[16177] = 8'h1b ;
            rom[16178] = 8'hdf ;
            rom[16179] = 8'hf2 ;
            rom[16180] = 8'h15 ;
            rom[16181] = 8'hfa ;
            rom[16182] = 8'hf9 ;
            rom[16183] = 8'h16 ;
            rom[16184] = 8'hf3 ;
            rom[16185] = 8'hef ;
            rom[16186] = 8'h1c ;
            rom[16187] = 8'h0f ;
            rom[16188] = 8'hff ;
            rom[16189] = 8'hde ;
            rom[16190] = 8'h16 ;
            rom[16191] = 8'hf7 ;
            rom[16192] = 8'h1c ;
            rom[16193] = 8'h04 ;
            rom[16194] = 8'he8 ;
            rom[16195] = 8'he9 ;
            rom[16196] = 8'h09 ;
            rom[16197] = 8'h0b ;
            rom[16198] = 8'h01 ;
            rom[16199] = 8'hd2 ;
            rom[16200] = 8'hff ;
            rom[16201] = 8'hfd ;
            rom[16202] = 8'h1c ;
            rom[16203] = 8'h28 ;
            rom[16204] = 8'h00 ;
            rom[16205] = 8'h04 ;
            rom[16206] = 8'hf9 ;
            rom[16207] = 8'hde ;
            rom[16208] = 8'h0c ;
            rom[16209] = 8'h00 ;
            rom[16210] = 8'hf0 ;
            rom[16211] = 8'hf7 ;
            rom[16212] = 8'hdf ;
            rom[16213] = 8'hd8 ;
            rom[16214] = 8'h0a ;
            rom[16215] = 8'hf6 ;
            rom[16216] = 8'h00 ;
            rom[16217] = 8'he7 ;
            rom[16218] = 8'h25 ;
            rom[16219] = 8'h08 ;
            rom[16220] = 8'hf9 ;
            rom[16221] = 8'he9 ;
            rom[16222] = 8'h07 ;
            rom[16223] = 8'h0f ;
            rom[16224] = 8'h13 ;
            rom[16225] = 8'h03 ;
            rom[16226] = 8'hfd ;
            rom[16227] = 8'hde ;
            rom[16228] = 8'h25 ;
            rom[16229] = 8'h2e ;
            rom[16230] = 8'he4 ;
            rom[16231] = 8'hdd ;
            rom[16232] = 8'h02 ;
            rom[16233] = 8'hf3 ;
            rom[16234] = 8'hfa ;
            rom[16235] = 8'h16 ;
            rom[16236] = 8'hec ;
            rom[16237] = 8'he9 ;
            rom[16238] = 8'he8 ;
            rom[16239] = 8'h0b ;
            rom[16240] = 8'he7 ;
            rom[16241] = 8'he1 ;
            rom[16242] = 8'h06 ;
            rom[16243] = 8'h00 ;
            rom[16244] = 8'hc5 ;
            rom[16245] = 8'he5 ;
            rom[16246] = 8'h23 ;
            rom[16247] = 8'h05 ;
            rom[16248] = 8'h02 ;
            rom[16249] = 8'h00 ;
            rom[16250] = 8'hfa ;
            rom[16251] = 8'h02 ;
            rom[16252] = 8'hee ;
            rom[16253] = 8'h02 ;
            rom[16254] = 8'h01 ;
            rom[16255] = 8'h02 ;
            rom[16256] = 8'h05 ;
            rom[16257] = 8'hfd ;
            rom[16258] = 8'he5 ;
            rom[16259] = 8'hf2 ;
            rom[16260] = 8'hff ;
            rom[16261] = 8'he5 ;
            rom[16262] = 8'hfb ;
            rom[16263] = 8'hfc ;
            rom[16264] = 8'hea ;
            rom[16265] = 8'h0b ;
            rom[16266] = 8'hff ;
            rom[16267] = 8'h28 ;
            rom[16268] = 8'hf1 ;
            rom[16269] = 8'he8 ;
            rom[16270] = 8'hfa ;
            rom[16271] = 8'hf2 ;
            rom[16272] = 8'h0b ;
            rom[16273] = 8'hf4 ;
            rom[16274] = 8'h09 ;
            rom[16275] = 8'h0e ;
            rom[16276] = 8'hff ;
            rom[16277] = 8'h22 ;
            rom[16278] = 8'hf6 ;
            rom[16279] = 8'hf3 ;
            rom[16280] = 8'hf2 ;
            rom[16281] = 8'hf0 ;
            rom[16282] = 8'h0a ;
            rom[16283] = 8'he4 ;
            rom[16284] = 8'he9 ;
            rom[16285] = 8'h08 ;
            rom[16286] = 8'h0c ;
            rom[16287] = 8'he5 ;
            rom[16288] = 8'he9 ;
            rom[16289] = 8'h0b ;
            rom[16290] = 8'hf7 ;
            rom[16291] = 8'hef ;
            rom[16292] = 8'hfb ;
            rom[16293] = 8'h22 ;
            rom[16294] = 8'hf2 ;
            rom[16295] = 8'h09 ;
            rom[16296] = 8'h0b ;
            rom[16297] = 8'h0b ;
            rom[16298] = 8'h1f ;
            rom[16299] = 8'hf4 ;
            rom[16300] = 8'hfe ;
            rom[16301] = 8'h10 ;
            rom[16302] = 8'h05 ;
            rom[16303] = 8'heb ;
            rom[16304] = 8'he0 ;
            rom[16305] = 8'hee ;
            rom[16306] = 8'he9 ;
            rom[16307] = 8'he3 ;
            rom[16308] = 8'hf2 ;
            rom[16309] = 8'h1b ;
            rom[16310] = 8'hf7 ;
            rom[16311] = 8'h25 ;
            rom[16312] = 8'hf5 ;
            rom[16313] = 8'h1b ;
            rom[16314] = 8'h14 ;
            rom[16315] = 8'h1e ;
            rom[16316] = 8'hfd ;
            rom[16317] = 8'hd2 ;
            rom[16318] = 8'hef ;
            rom[16319] = 8'h1e ;
            rom[16320] = 8'hee ;
            rom[16321] = 8'hff ;
            rom[16322] = 8'hf2 ;
            rom[16323] = 8'h12 ;
            rom[16324] = 8'h02 ;
            rom[16325] = 8'h00 ;
            rom[16326] = 8'hf7 ;
            rom[16327] = 8'h0e ;
            rom[16328] = 8'h00 ;
            rom[16329] = 8'hf9 ;
            rom[16330] = 8'hf9 ;
            rom[16331] = 8'h00 ;
            rom[16332] = 8'h0d ;
            rom[16333] = 8'hee ;
            rom[16334] = 8'h1d ;
            rom[16335] = 8'hd3 ;
            rom[16336] = 8'hf6 ;
            rom[16337] = 8'h08 ;
            rom[16338] = 8'h0f ;
            rom[16339] = 8'hf7 ;
            rom[16340] = 8'he6 ;
            rom[16341] = 8'hfd ;
            rom[16342] = 8'h0e ;
            rom[16343] = 8'h0b ;
            rom[16344] = 8'hfb ;
            rom[16345] = 8'h1b ;
            rom[16346] = 8'h09 ;
            rom[16347] = 8'he9 ;
            rom[16348] = 8'h1a ;
            rom[16349] = 8'he5 ;
            rom[16350] = 8'hfb ;
            rom[16351] = 8'h0d ;
            rom[16352] = 8'hf2 ;
            rom[16353] = 8'h02 ;
            rom[16354] = 8'he3 ;
            rom[16355] = 8'heb ;
            rom[16356] = 8'h24 ;
            rom[16357] = 8'h25 ;
            rom[16358] = 8'h19 ;
            rom[16359] = 8'hf2 ;
            rom[16360] = 8'hfc ;
            rom[16361] = 8'hfb ;
            rom[16362] = 8'h14 ;
            rom[16363] = 8'h19 ;
            rom[16364] = 8'h04 ;
            rom[16365] = 8'hf2 ;
            rom[16366] = 8'h28 ;
            rom[16367] = 8'h03 ;
            rom[16368] = 8'hfc ;
            rom[16369] = 8'hfe ;
            rom[16370] = 8'h05 ;
            rom[16371] = 8'h05 ;
            rom[16372] = 8'hff ;
            rom[16373] = 8'hfb ;
            rom[16374] = 8'h0b ;
            rom[16375] = 8'h00 ;
            rom[16376] = 8'h22 ;
            rom[16377] = 8'hf7 ;
            rom[16378] = 8'h21 ;
            rom[16379] = 8'hfa ;
            rom[16380] = 8'h13 ;
            rom[16381] = 8'h0c ;
            rom[16382] = 8'hf4 ;
            rom[16383] = 8'hdb ;
            rom[16384] = 8'h21 ;
            rom[16385] = 8'h02 ;
            rom[16386] = 8'hdc ;
            rom[16387] = 8'hec ;
            rom[16388] = 8'h15 ;
            rom[16389] = 8'hf2 ;
            rom[16390] = 8'h13 ;
            rom[16391] = 8'hd5 ;
            rom[16392] = 8'hf8 ;
            rom[16393] = 8'h12 ;
            rom[16394] = 8'hee ;
            rom[16395] = 8'hf0 ;
            rom[16396] = 8'hfb ;
            rom[16397] = 8'h23 ;
            rom[16398] = 8'h0d ;
            rom[16399] = 8'hdb ;
            rom[16400] = 8'h07 ;
            rom[16401] = 8'h07 ;
            rom[16402] = 8'hf7 ;
            rom[16403] = 8'hf3 ;
            rom[16404] = 8'hea ;
            rom[16405] = 8'h0d ;
            rom[16406] = 8'he9 ;
            rom[16407] = 8'h04 ;
            rom[16408] = 8'h06 ;
            rom[16409] = 8'h00 ;
            rom[16410] = 8'h01 ;
            rom[16411] = 8'hff ;
            rom[16412] = 8'hfa ;
            rom[16413] = 8'hff ;
            rom[16414] = 8'hed ;
            rom[16415] = 8'hf5 ;
            rom[16416] = 8'he8 ;
            rom[16417] = 8'hee ;
            rom[16418] = 8'hf5 ;
            rom[16419] = 8'h04 ;
            rom[16420] = 8'h0e ;
            rom[16421] = 8'h0e ;
            rom[16422] = 8'hcc ;
            rom[16423] = 8'hdd ;
            rom[16424] = 8'h1f ;
            rom[16425] = 8'h07 ;
            rom[16426] = 8'h08 ;
            rom[16427] = 8'he8 ;
            rom[16428] = 8'hfd ;
            rom[16429] = 8'hf7 ;
            rom[16430] = 8'h13 ;
            rom[16431] = 8'hfc ;
            rom[16432] = 8'he9 ;
            rom[16433] = 8'h16 ;
            rom[16434] = 8'h0b ;
            rom[16435] = 8'hf1 ;
            rom[16436] = 8'hf6 ;
            rom[16437] = 8'hfc ;
            rom[16438] = 8'he6 ;
            rom[16439] = 8'hfd ;
            rom[16440] = 8'hf4 ;
            rom[16441] = 8'hf8 ;
            rom[16442] = 8'h04 ;
            rom[16443] = 8'hfb ;
            rom[16444] = 8'hdd ;
            rom[16445] = 8'h00 ;
            rom[16446] = 8'hda ;
            rom[16447] = 8'h03 ;
            rom[16448] = 8'h10 ;
            rom[16449] = 8'he2 ;
            rom[16450] = 8'h34 ;
            rom[16451] = 8'hf5 ;
            rom[16452] = 8'h19 ;
            rom[16453] = 8'h01 ;
            rom[16454] = 8'h1e ;
            rom[16455] = 8'h11 ;
            rom[16456] = 8'hda ;
            rom[16457] = 8'h25 ;
            rom[16458] = 8'he3 ;
            rom[16459] = 8'he3 ;
            rom[16460] = 8'h0f ;
            rom[16461] = 8'h1b ;
            rom[16462] = 8'hfc ;
            rom[16463] = 8'hdd ;
            rom[16464] = 8'hf6 ;
            rom[16465] = 8'h0b ;
            rom[16466] = 8'h2b ;
            rom[16467] = 8'h0c ;
            rom[16468] = 8'hef ;
            rom[16469] = 8'hec ;
            rom[16470] = 8'hfb ;
            rom[16471] = 8'h26 ;
            rom[16472] = 8'hf3 ;
            rom[16473] = 8'hfa ;
            rom[16474] = 8'hfc ;
            rom[16475] = 8'h11 ;
            rom[16476] = 8'hf9 ;
            rom[16477] = 8'heb ;
            rom[16478] = 8'h14 ;
            rom[16479] = 8'hfa ;
            rom[16480] = 8'h08 ;
            rom[16481] = 8'hf4 ;
            rom[16482] = 8'hfa ;
            rom[16483] = 8'h24 ;
            rom[16484] = 8'hf0 ;
            rom[16485] = 8'hdf ;
            rom[16486] = 8'heb ;
            rom[16487] = 8'hfe ;
            rom[16488] = 8'hf0 ;
            rom[16489] = 8'h15 ;
            rom[16490] = 8'h29 ;
            rom[16491] = 8'hf1 ;
            rom[16492] = 8'h10 ;
            rom[16493] = 8'hf7 ;
            rom[16494] = 8'hf5 ;
            rom[16495] = 8'h11 ;
            rom[16496] = 8'he9 ;
            rom[16497] = 8'hfc ;
            rom[16498] = 8'hfe ;
            rom[16499] = 8'hed ;
            rom[16500] = 8'hf5 ;
            rom[16501] = 8'h16 ;
            rom[16502] = 8'h16 ;
            rom[16503] = 8'h01 ;
            rom[16504] = 8'hec ;
            rom[16505] = 8'h07 ;
            rom[16506] = 8'hf2 ;
            rom[16507] = 8'hdd ;
            rom[16508] = 8'h06 ;
            rom[16509] = 8'h16 ;
            rom[16510] = 8'hfc ;
            rom[16511] = 8'h22 ;
            rom[16512] = 8'h04 ;
            rom[16513] = 8'hf8 ;
            rom[16514] = 8'h14 ;
            rom[16515] = 8'h1a ;
            rom[16516] = 8'hf9 ;
            rom[16517] = 8'he1 ;
            rom[16518] = 8'hcd ;
            rom[16519] = 8'h12 ;
            rom[16520] = 8'h0a ;
            rom[16521] = 8'he8 ;
            rom[16522] = 8'h0a ;
            rom[16523] = 8'h13 ;
            rom[16524] = 8'h06 ;
            rom[16525] = 8'hf7 ;
            rom[16526] = 8'h00 ;
            rom[16527] = 8'hd4 ;
            rom[16528] = 8'he6 ;
            rom[16529] = 8'hfa ;
            rom[16530] = 8'h11 ;
            rom[16531] = 8'h06 ;
            rom[16532] = 8'h08 ;
            rom[16533] = 8'h21 ;
            rom[16534] = 8'hee ;
            rom[16535] = 8'h02 ;
            rom[16536] = 8'h3d ;
            rom[16537] = 8'h1a ;
            rom[16538] = 8'h04 ;
            rom[16539] = 8'h12 ;
            rom[16540] = 8'hff ;
            rom[16541] = 8'h11 ;
            rom[16542] = 8'hff ;
            rom[16543] = 8'hee ;
            rom[16544] = 8'h05 ;
            rom[16545] = 8'he4 ;
            rom[16546] = 8'hf4 ;
            rom[16547] = 8'hf6 ;
            rom[16548] = 8'h11 ;
            rom[16549] = 8'h09 ;
            rom[16550] = 8'hfa ;
            rom[16551] = 8'hb5 ;
            rom[16552] = 8'h00 ;
            rom[16553] = 8'hec ;
            rom[16554] = 8'hf6 ;
            rom[16555] = 8'hf3 ;
            rom[16556] = 8'hf2 ;
            rom[16557] = 8'h05 ;
            rom[16558] = 8'hf4 ;
            rom[16559] = 8'he4 ;
            rom[16560] = 8'h08 ;
            rom[16561] = 8'hf9 ;
            rom[16562] = 8'h06 ;
            rom[16563] = 8'hf2 ;
            rom[16564] = 8'h04 ;
            rom[16565] = 8'h25 ;
            rom[16566] = 8'hea ;
            rom[16567] = 8'hf2 ;
            rom[16568] = 8'h09 ;
            rom[16569] = 8'h0a ;
            rom[16570] = 8'h04 ;
            rom[16571] = 8'hf0 ;
            rom[16572] = 8'h21 ;
            rom[16573] = 8'hf2 ;
            rom[16574] = 8'h2d ;
            rom[16575] = 8'he8 ;
            rom[16576] = 8'hfa ;
            rom[16577] = 8'h0f ;
            rom[16578] = 8'hf9 ;
            rom[16579] = 8'hf6 ;
            rom[16580] = 8'h01 ;
            rom[16581] = 8'hfe ;
            rom[16582] = 8'hfb ;
            rom[16583] = 8'h0d ;
            rom[16584] = 8'h0b ;
            rom[16585] = 8'hf4 ;
            rom[16586] = 8'h0a ;
            rom[16587] = 8'hf9 ;
            rom[16588] = 8'hfc ;
            rom[16589] = 8'hf6 ;
            rom[16590] = 8'h17 ;
            rom[16591] = 8'hf4 ;
            rom[16592] = 8'h09 ;
            rom[16593] = 8'hdb ;
            rom[16594] = 8'h02 ;
            rom[16595] = 8'hf1 ;
            rom[16596] = 8'h0a ;
            rom[16597] = 8'hc8 ;
            rom[16598] = 8'he2 ;
            rom[16599] = 8'hd9 ;
            rom[16600] = 8'h0e ;
            rom[16601] = 8'hfe ;
            rom[16602] = 8'h28 ;
            rom[16603] = 8'hfe ;
            rom[16604] = 8'h17 ;
            rom[16605] = 8'h00 ;
            rom[16606] = 8'hf6 ;
            rom[16607] = 8'hdc ;
            rom[16608] = 8'heb ;
            rom[16609] = 8'h1b ;
            rom[16610] = 8'hf8 ;
            rom[16611] = 8'hf2 ;
            rom[16612] = 8'h01 ;
            rom[16613] = 8'he3 ;
            rom[16614] = 8'hec ;
            rom[16615] = 8'hfb ;
            rom[16616] = 8'h02 ;
            rom[16617] = 8'h0a ;
            rom[16618] = 8'h24 ;
            rom[16619] = 8'he4 ;
            rom[16620] = 8'hfc ;
            rom[16621] = 8'he7 ;
            rom[16622] = 8'hdf ;
            rom[16623] = 8'hf0 ;
            rom[16624] = 8'h1d ;
            rom[16625] = 8'hea ;
            rom[16626] = 8'h05 ;
            rom[16627] = 8'hed ;
            rom[16628] = 8'hf3 ;
            rom[16629] = 8'h16 ;
            rom[16630] = 8'h2a ;
            rom[16631] = 8'hf2 ;
            rom[16632] = 8'h20 ;
            rom[16633] = 8'hfd ;
            rom[16634] = 8'h0e ;
            rom[16635] = 8'hfd ;
            rom[16636] = 8'h0c ;
            rom[16637] = 8'hf7 ;
            rom[16638] = 8'he1 ;
            rom[16639] = 8'hff ;
            rom[16640] = 8'h24 ;
            rom[16641] = 8'h14 ;
            rom[16642] = 8'hf9 ;
            rom[16643] = 8'h0c ;
            rom[16644] = 8'hf1 ;
            rom[16645] = 8'h05 ;
            rom[16646] = 8'h20 ;
            rom[16647] = 8'h2e ;
            rom[16648] = 8'h04 ;
            rom[16649] = 8'h2a ;
            rom[16650] = 8'hf7 ;
            rom[16651] = 8'heb ;
            rom[16652] = 8'h00 ;
            rom[16653] = 8'h03 ;
            rom[16654] = 8'h04 ;
            rom[16655] = 8'h0e ;
            rom[16656] = 8'hb5 ;
            rom[16657] = 8'hd3 ;
            rom[16658] = 8'h0d ;
            rom[16659] = 8'h15 ;
            rom[16660] = 8'hd7 ;
            rom[16661] = 8'he7 ;
            rom[16662] = 8'hea ;
            rom[16663] = 8'h04 ;
            rom[16664] = 8'h09 ;
            rom[16665] = 8'h07 ;
            rom[16666] = 8'hf5 ;
            rom[16667] = 8'hfb ;
            rom[16668] = 8'hf5 ;
            rom[16669] = 8'he1 ;
            rom[16670] = 8'hf8 ;
            rom[16671] = 8'hfc ;
            rom[16672] = 8'hf8 ;
            rom[16673] = 8'he1 ;
            rom[16674] = 8'he8 ;
            rom[16675] = 8'hec ;
            rom[16676] = 8'hec ;
            rom[16677] = 8'hff ;
            rom[16678] = 8'hd5 ;
            rom[16679] = 8'hfe ;
            rom[16680] = 8'hfd ;
            rom[16681] = 8'h2f ;
            rom[16682] = 8'he1 ;
            rom[16683] = 8'hfd ;
            rom[16684] = 8'hdb ;
            rom[16685] = 8'hf3 ;
            rom[16686] = 8'hde ;
            rom[16687] = 8'hf6 ;
            rom[16688] = 8'hea ;
            rom[16689] = 8'h0b ;
            rom[16690] = 8'hf4 ;
            rom[16691] = 8'hf7 ;
            rom[16692] = 8'h06 ;
            rom[16693] = 8'h0d ;
            rom[16694] = 8'hf7 ;
            rom[16695] = 8'hdf ;
            rom[16696] = 8'h12 ;
            rom[16697] = 8'hff ;
            rom[16698] = 8'h11 ;
            rom[16699] = 8'hfe ;
            rom[16700] = 8'h0c ;
            rom[16701] = 8'hfe ;
            rom[16702] = 8'he9 ;
            rom[16703] = 8'hf9 ;
            rom[16704] = 8'h0b ;
            rom[16705] = 8'hd0 ;
            rom[16706] = 8'hf5 ;
            rom[16707] = 8'h07 ;
            rom[16708] = 8'hec ;
            rom[16709] = 8'h10 ;
            rom[16710] = 8'h00 ;
            rom[16711] = 8'hf4 ;
            rom[16712] = 8'h0d ;
            rom[16713] = 8'h1b ;
            rom[16714] = 8'h30 ;
            rom[16715] = 8'h10 ;
            rom[16716] = 8'hf2 ;
            rom[16717] = 8'h04 ;
            rom[16718] = 8'he7 ;
            rom[16719] = 8'hff ;
            rom[16720] = 8'hf9 ;
            rom[16721] = 8'heb ;
            rom[16722] = 8'hf7 ;
            rom[16723] = 8'he7 ;
            rom[16724] = 8'hf9 ;
            rom[16725] = 8'h0a ;
            rom[16726] = 8'h19 ;
            rom[16727] = 8'h0a ;
            rom[16728] = 8'hf9 ;
            rom[16729] = 8'hdd ;
            rom[16730] = 8'h1d ;
            rom[16731] = 8'hed ;
            rom[16732] = 8'h01 ;
            rom[16733] = 8'hd9 ;
            rom[16734] = 8'ha8 ;
            rom[16735] = 8'h11 ;
            rom[16736] = 8'heb ;
            rom[16737] = 8'h10 ;
            rom[16738] = 8'he8 ;
            rom[16739] = 8'he7 ;
            rom[16740] = 8'h02 ;
            rom[16741] = 8'he4 ;
            rom[16742] = 8'h16 ;
            rom[16743] = 8'h16 ;
            rom[16744] = 8'hdf ;
            rom[16745] = 8'hf7 ;
            rom[16746] = 8'hd5 ;
            rom[16747] = 8'h08 ;
            rom[16748] = 8'hf4 ;
            rom[16749] = 8'hfe ;
            rom[16750] = 8'h13 ;
            rom[16751] = 8'hfb ;
            rom[16752] = 8'h04 ;
            rom[16753] = 8'hf7 ;
            rom[16754] = 8'heb ;
            rom[16755] = 8'hdc ;
            rom[16756] = 8'h10 ;
            rom[16757] = 8'h07 ;
            rom[16758] = 8'hea ;
            rom[16759] = 8'h05 ;
            rom[16760] = 8'h0f ;
            rom[16761] = 8'h06 ;
            rom[16762] = 8'h0e ;
            rom[16763] = 8'heb ;
            rom[16764] = 8'h0e ;
            rom[16765] = 8'h0c ;
            rom[16766] = 8'h18 ;
            rom[16767] = 8'hde ;
            rom[16768] = 8'hdb ;
            rom[16769] = 8'h16 ;
            rom[16770] = 8'hfc ;
            rom[16771] = 8'h19 ;
            rom[16772] = 8'h03 ;
            rom[16773] = 8'hda ;
            rom[16774] = 8'hfc ;
            rom[16775] = 8'h13 ;
            rom[16776] = 8'h03 ;
            rom[16777] = 8'hfb ;
            rom[16778] = 8'h0f ;
            rom[16779] = 8'h0e ;
            rom[16780] = 8'hd3 ;
            rom[16781] = 8'h04 ;
            rom[16782] = 8'h05 ;
            rom[16783] = 8'h0d ;
            rom[16784] = 8'hf5 ;
            rom[16785] = 8'h16 ;
            rom[16786] = 8'he5 ;
            rom[16787] = 8'h19 ;
            rom[16788] = 8'h0e ;
            rom[16789] = 8'h17 ;
            rom[16790] = 8'hd3 ;
            rom[16791] = 8'hfb ;
            rom[16792] = 8'h03 ;
            rom[16793] = 8'hf9 ;
            rom[16794] = 8'h03 ;
            rom[16795] = 8'h14 ;
            rom[16796] = 8'he8 ;
            rom[16797] = 8'h23 ;
            rom[16798] = 8'h03 ;
            rom[16799] = 8'hf5 ;
            rom[16800] = 8'h03 ;
            rom[16801] = 8'hcb ;
            rom[16802] = 8'h13 ;
            rom[16803] = 8'h05 ;
            rom[16804] = 8'h12 ;
            rom[16805] = 8'he5 ;
            rom[16806] = 8'hf0 ;
            rom[16807] = 8'he2 ;
            rom[16808] = 8'h08 ;
            rom[16809] = 8'h06 ;
            rom[16810] = 8'h04 ;
            rom[16811] = 8'hfd ;
            rom[16812] = 8'he9 ;
            rom[16813] = 8'hdc ;
            rom[16814] = 8'hf2 ;
            rom[16815] = 8'he6 ;
            rom[16816] = 8'h12 ;
            rom[16817] = 8'hfb ;
            rom[16818] = 8'hbb ;
            rom[16819] = 8'he8 ;
            rom[16820] = 8'h0a ;
            rom[16821] = 8'h0f ;
            rom[16822] = 8'h11 ;
            rom[16823] = 8'hdd ;
            rom[16824] = 8'hfd ;
            rom[16825] = 8'h25 ;
            rom[16826] = 8'h13 ;
            rom[16827] = 8'hea ;
            rom[16828] = 8'hfe ;
            rom[16829] = 8'hf8 ;
            rom[16830] = 8'h12 ;
            rom[16831] = 8'hfb ;
            rom[16832] = 8'hff ;
            rom[16833] = 8'h30 ;
            rom[16834] = 8'hd0 ;
            rom[16835] = 8'h11 ;
            rom[16836] = 8'hf4 ;
            rom[16837] = 8'hf6 ;
            rom[16838] = 8'hf5 ;
            rom[16839] = 8'h44 ;
            rom[16840] = 8'h18 ;
            rom[16841] = 8'h1e ;
            rom[16842] = 8'hfe ;
            rom[16843] = 8'hf4 ;
            rom[16844] = 8'hf1 ;
            rom[16845] = 8'he6 ;
            rom[16846] = 8'h27 ;
            rom[16847] = 8'hf3 ;
            rom[16848] = 8'h01 ;
            rom[16849] = 8'hd9 ;
            rom[16850] = 8'h08 ;
            rom[16851] = 8'h11 ;
            rom[16852] = 8'h03 ;
            rom[16853] = 8'hfa ;
            rom[16854] = 8'heb ;
            rom[16855] = 8'h0a ;
            rom[16856] = 8'hfd ;
            rom[16857] = 8'hfa ;
            rom[16858] = 8'h08 ;
            rom[16859] = 8'hed ;
            rom[16860] = 8'hfc ;
            rom[16861] = 8'h18 ;
            rom[16862] = 8'hd3 ;
            rom[16863] = 8'he5 ;
            rom[16864] = 8'he9 ;
            rom[16865] = 8'hd1 ;
            rom[16866] = 8'hde ;
            rom[16867] = 8'h00 ;
            rom[16868] = 8'h17 ;
            rom[16869] = 8'hda ;
            rom[16870] = 8'hfd ;
            rom[16871] = 8'hd8 ;
            rom[16872] = 8'h02 ;
            rom[16873] = 8'h28 ;
            rom[16874] = 8'hdf ;
            rom[16875] = 8'h0c ;
            rom[16876] = 8'hc6 ;
            rom[16877] = 8'h12 ;
            rom[16878] = 8'he1 ;
            rom[16879] = 8'he8 ;
            rom[16880] = 8'h11 ;
            rom[16881] = 8'hdf ;
            rom[16882] = 8'h1b ;
            rom[16883] = 8'hc4 ;
            rom[16884] = 8'h0c ;
            rom[16885] = 8'h18 ;
            rom[16886] = 8'h07 ;
            rom[16887] = 8'hef ;
            rom[16888] = 8'hdb ;
            rom[16889] = 8'hf5 ;
            rom[16890] = 8'h1a ;
            rom[16891] = 8'h08 ;
            rom[16892] = 8'h0b ;
            rom[16893] = 8'hed ;
            rom[16894] = 8'h13 ;
            rom[16895] = 8'hed ;
            rom[16896] = 8'h09 ;
            rom[16897] = 8'hde ;
            rom[16898] = 8'h0d ;
            rom[16899] = 8'hec ;
            rom[16900] = 8'hce ;
            rom[16901] = 8'h02 ;
            rom[16902] = 8'h0f ;
            rom[16903] = 8'h0c ;
            rom[16904] = 8'he5 ;
            rom[16905] = 8'h0d ;
            rom[16906] = 8'h02 ;
            rom[16907] = 8'hfc ;
            rom[16908] = 8'h0a ;
            rom[16909] = 8'h05 ;
            rom[16910] = 8'h1b ;
            rom[16911] = 8'h06 ;
            rom[16912] = 8'hbd ;
            rom[16913] = 8'hfb ;
            rom[16914] = 8'h1f ;
            rom[16915] = 8'hfc ;
            rom[16916] = 8'hd6 ;
            rom[16917] = 8'he7 ;
            rom[16918] = 8'hf9 ;
            rom[16919] = 8'h08 ;
            rom[16920] = 8'hf8 ;
            rom[16921] = 8'hd2 ;
            rom[16922] = 8'h02 ;
            rom[16923] = 8'hf6 ;
            rom[16924] = 8'hf5 ;
            rom[16925] = 8'hc4 ;
            rom[16926] = 8'h08 ;
            rom[16927] = 8'hdc ;
            rom[16928] = 8'h06 ;
            rom[16929] = 8'hc9 ;
            rom[16930] = 8'hff ;
            rom[16931] = 8'he3 ;
            rom[16932] = 8'h04 ;
            rom[16933] = 8'he5 ;
            rom[16934] = 8'h10 ;
            rom[16935] = 8'hef ;
            rom[16936] = 8'hea ;
            rom[16937] = 8'h2c ;
            rom[16938] = 8'h17 ;
            rom[16939] = 8'hfa ;
            rom[16940] = 8'h23 ;
            rom[16941] = 8'h1b ;
            rom[16942] = 8'h0f ;
            rom[16943] = 8'hec ;
            rom[16944] = 8'hff ;
            rom[16945] = 8'hf9 ;
            rom[16946] = 8'hd2 ;
            rom[16947] = 8'hf9 ;
            rom[16948] = 8'h0a ;
            rom[16949] = 8'h01 ;
            rom[16950] = 8'hf9 ;
            rom[16951] = 8'hdf ;
            rom[16952] = 8'h11 ;
            rom[16953] = 8'h05 ;
            rom[16954] = 8'h0c ;
            rom[16955] = 8'hfc ;
            rom[16956] = 8'h01 ;
            rom[16957] = 8'hfa ;
            rom[16958] = 8'h08 ;
            rom[16959] = 8'h1a ;
            rom[16960] = 8'h13 ;
            rom[16961] = 8'he7 ;
            rom[16962] = 8'h06 ;
            rom[16963] = 8'hfc ;
            rom[16964] = 8'hf4 ;
            rom[16965] = 8'hfb ;
            rom[16966] = 8'h0c ;
            rom[16967] = 8'h06 ;
            rom[16968] = 8'hff ;
            rom[16969] = 8'h00 ;
            rom[16970] = 8'h00 ;
            rom[16971] = 8'h01 ;
            rom[16972] = 8'h16 ;
            rom[16973] = 8'h0c ;
            rom[16974] = 8'h0f ;
            rom[16975] = 8'hea ;
            rom[16976] = 8'hd7 ;
            rom[16977] = 8'h07 ;
            rom[16978] = 8'h0b ;
            rom[16979] = 8'h04 ;
            rom[16980] = 8'h06 ;
            rom[16981] = 8'hdc ;
            rom[16982] = 8'h0e ;
            rom[16983] = 8'h1e ;
            rom[16984] = 8'h0b ;
            rom[16985] = 8'h03 ;
            rom[16986] = 8'hf3 ;
            rom[16987] = 8'h06 ;
            rom[16988] = 8'h07 ;
            rom[16989] = 8'hf3 ;
            rom[16990] = 8'h10 ;
            rom[16991] = 8'hfb ;
            rom[16992] = 8'hfa ;
            rom[16993] = 8'hf5 ;
            rom[16994] = 8'hf7 ;
            rom[16995] = 8'hfb ;
            rom[16996] = 8'hff ;
            rom[16997] = 8'hfc ;
            rom[16998] = 8'hfa ;
            rom[16999] = 8'hf7 ;
            rom[17000] = 8'hfa ;
            rom[17001] = 8'h26 ;
            rom[17002] = 8'h03 ;
            rom[17003] = 8'hfe ;
            rom[17004] = 8'h16 ;
            rom[17005] = 8'h0e ;
            rom[17006] = 8'h0c ;
            rom[17007] = 8'hfa ;
            rom[17008] = 8'hda ;
            rom[17009] = 8'hff ;
            rom[17010] = 8'hd3 ;
            rom[17011] = 8'hf0 ;
            rom[17012] = 8'h18 ;
            rom[17013] = 8'h14 ;
            rom[17014] = 8'h13 ;
            rom[17015] = 8'he6 ;
            rom[17016] = 8'h11 ;
            rom[17017] = 8'h15 ;
            rom[17018] = 8'hf6 ;
            rom[17019] = 8'hed ;
            rom[17020] = 8'h23 ;
            rom[17021] = 8'h04 ;
            rom[17022] = 8'hfc ;
            rom[17023] = 8'h22 ;
            rom[17024] = 8'hf5 ;
            rom[17025] = 8'hdb ;
            rom[17026] = 8'h1e ;
            rom[17027] = 8'h07 ;
            rom[17028] = 8'hfe ;
            rom[17029] = 8'h04 ;
            rom[17030] = 8'h0c ;
            rom[17031] = 8'h02 ;
            rom[17032] = 8'h07 ;
            rom[17033] = 8'hfd ;
            rom[17034] = 8'hfc ;
            rom[17035] = 8'h10 ;
            rom[17036] = 8'hfc ;
            rom[17037] = 8'hf4 ;
            rom[17038] = 8'h04 ;
            rom[17039] = 8'h17 ;
            rom[17040] = 8'hfc ;
            rom[17041] = 8'h10 ;
            rom[17042] = 8'h1a ;
            rom[17043] = 8'h21 ;
            rom[17044] = 8'h05 ;
            rom[17045] = 8'h0f ;
            rom[17046] = 8'hf9 ;
            rom[17047] = 8'hde ;
            rom[17048] = 8'h17 ;
            rom[17049] = 8'he5 ;
            rom[17050] = 8'hf5 ;
            rom[17051] = 8'hd2 ;
            rom[17052] = 8'hf0 ;
            rom[17053] = 8'hf2 ;
            rom[17054] = 8'he6 ;
            rom[17055] = 8'h04 ;
            rom[17056] = 8'he9 ;
            rom[17057] = 8'hf5 ;
            rom[17058] = 8'hf6 ;
            rom[17059] = 8'hef ;
            rom[17060] = 8'hf8 ;
            rom[17061] = 8'he8 ;
            rom[17062] = 8'h25 ;
            rom[17063] = 8'h06 ;
            rom[17064] = 8'heb ;
            rom[17065] = 8'h02 ;
            rom[17066] = 8'hf8 ;
            rom[17067] = 8'hf0 ;
            rom[17068] = 8'h0a ;
            rom[17069] = 8'hf9 ;
            rom[17070] = 8'h29 ;
            rom[17071] = 8'h1a ;
            rom[17072] = 8'hf3 ;
            rom[17073] = 8'hf6 ;
            rom[17074] = 8'h13 ;
            rom[17075] = 8'hdd ;
            rom[17076] = 8'h1e ;
            rom[17077] = 8'he9 ;
            rom[17078] = 8'hdc ;
            rom[17079] = 8'h11 ;
            rom[17080] = 8'h0a ;
            rom[17081] = 8'h00 ;
            rom[17082] = 8'h12 ;
            rom[17083] = 8'h2d ;
            rom[17084] = 8'h09 ;
            rom[17085] = 8'h16 ;
            rom[17086] = 8'h0d ;
            rom[17087] = 8'h06 ;
            rom[17088] = 8'h16 ;
            rom[17089] = 8'h05 ;
            rom[17090] = 8'h16 ;
            rom[17091] = 8'hd9 ;
            rom[17092] = 8'hda ;
            rom[17093] = 8'hef ;
            rom[17094] = 8'h04 ;
            rom[17095] = 8'hfc ;
            rom[17096] = 8'heb ;
            rom[17097] = 8'h21 ;
            rom[17098] = 8'hff ;
            rom[17099] = 8'h29 ;
            rom[17100] = 8'h00 ;
            rom[17101] = 8'h11 ;
            rom[17102] = 8'h2c ;
            rom[17103] = 8'h14 ;
            rom[17104] = 8'hf4 ;
            rom[17105] = 8'hcf ;
            rom[17106] = 8'h17 ;
            rom[17107] = 8'hec ;
            rom[17108] = 8'hed ;
            rom[17109] = 8'h14 ;
            rom[17110] = 8'hce ;
            rom[17111] = 8'hfd ;
            rom[17112] = 8'h2c ;
            rom[17113] = 8'hfa ;
            rom[17114] = 8'h1b ;
            rom[17115] = 8'h0e ;
            rom[17116] = 8'h2a ;
            rom[17117] = 8'hd7 ;
            rom[17118] = 8'h17 ;
            rom[17119] = 8'heb ;
            rom[17120] = 8'h13 ;
            rom[17121] = 8'hec ;
            rom[17122] = 8'h06 ;
            rom[17123] = 8'h03 ;
            rom[17124] = 8'hdd ;
            rom[17125] = 8'h0a ;
            rom[17126] = 8'hf4 ;
            rom[17127] = 8'h07 ;
            rom[17128] = 8'hf5 ;
            rom[17129] = 8'hfc ;
            rom[17130] = 8'h02 ;
            rom[17131] = 8'hfe ;
            rom[17132] = 8'hf9 ;
            rom[17133] = 8'hd5 ;
            rom[17134] = 8'he4 ;
            rom[17135] = 8'h04 ;
            rom[17136] = 8'he2 ;
            rom[17137] = 8'hda ;
            rom[17138] = 8'hda ;
            rom[17139] = 8'hf7 ;
            rom[17140] = 8'h1a ;
            rom[17141] = 8'h05 ;
            rom[17142] = 8'he7 ;
            rom[17143] = 8'h2f ;
            rom[17144] = 8'h1b ;
            rom[17145] = 8'h19 ;
            rom[17146] = 8'hfc ;
            rom[17147] = 8'he4 ;
            rom[17148] = 8'he7 ;
            rom[17149] = 8'h08 ;
            rom[17150] = 8'h15 ;
            rom[17151] = 8'h0d ;
            rom[17152] = 8'hfa ;
            rom[17153] = 8'h25 ;
            rom[17154] = 8'hfd ;
            rom[17155] = 8'heb ;
            rom[17156] = 8'h01 ;
            rom[17157] = 8'h08 ;
            rom[17158] = 8'hfa ;
            rom[17159] = 8'h0f ;
            rom[17160] = 8'he2 ;
            rom[17161] = 8'h20 ;
            rom[17162] = 8'h0a ;
            rom[17163] = 8'he7 ;
            rom[17164] = 8'he3 ;
            rom[17165] = 8'hf7 ;
            rom[17166] = 8'h0e ;
            rom[17167] = 8'h10 ;
            rom[17168] = 8'h02 ;
            rom[17169] = 8'h0f ;
            rom[17170] = 8'h03 ;
            rom[17171] = 8'h07 ;
            rom[17172] = 8'h07 ;
            rom[17173] = 8'h13 ;
            rom[17174] = 8'h0b ;
            rom[17175] = 8'h0a ;
            rom[17176] = 8'heb ;
            rom[17177] = 8'hf3 ;
            rom[17178] = 8'he0 ;
            rom[17179] = 8'h17 ;
            rom[17180] = 8'hf5 ;
            rom[17181] = 8'h1e ;
            rom[17182] = 8'h0a ;
            rom[17183] = 8'hdc ;
            rom[17184] = 8'h32 ;
            rom[17185] = 8'hd4 ;
            rom[17186] = 8'h0e ;
            rom[17187] = 8'h17 ;
            rom[17188] = 8'h0f ;
            rom[17189] = 8'hf9 ;
            rom[17190] = 8'hea ;
            rom[17191] = 8'he8 ;
            rom[17192] = 8'h0e ;
            rom[17193] = 8'h21 ;
            rom[17194] = 8'h0b ;
            rom[17195] = 8'h0f ;
            rom[17196] = 8'h11 ;
            rom[17197] = 8'h16 ;
            rom[17198] = 8'hf0 ;
            rom[17199] = 8'heb ;
            rom[17200] = 8'hee ;
            rom[17201] = 8'h04 ;
            rom[17202] = 8'hda ;
            rom[17203] = 8'he9 ;
            rom[17204] = 8'hfd ;
            rom[17205] = 8'h17 ;
            rom[17206] = 8'h07 ;
            rom[17207] = 8'hdb ;
            rom[17208] = 8'heb ;
            rom[17209] = 8'h1a ;
            rom[17210] = 8'hf3 ;
            rom[17211] = 8'h00 ;
            rom[17212] = 8'h09 ;
            rom[17213] = 8'hec ;
            rom[17214] = 8'h3c ;
            rom[17215] = 8'hff ;
            rom[17216] = 8'hf8 ;
            rom[17217] = 8'h04 ;
            rom[17218] = 8'hf1 ;
            rom[17219] = 8'he2 ;
            rom[17220] = 8'he9 ;
            rom[17221] = 8'h06 ;
            rom[17222] = 8'h2b ;
            rom[17223] = 8'he3 ;
            rom[17224] = 8'h06 ;
            rom[17225] = 8'h14 ;
            rom[17226] = 8'hff ;
            rom[17227] = 8'hd8 ;
            rom[17228] = 8'hfb ;
            rom[17229] = 8'h08 ;
            rom[17230] = 8'hf5 ;
            rom[17231] = 8'hf8 ;
            rom[17232] = 8'h07 ;
            rom[17233] = 8'hf3 ;
            rom[17234] = 8'h03 ;
            rom[17235] = 8'hd5 ;
            rom[17236] = 8'hdf ;
            rom[17237] = 8'hff ;
            rom[17238] = 8'h09 ;
            rom[17239] = 8'h0f ;
            rom[17240] = 8'hf3 ;
            rom[17241] = 8'hf3 ;
            rom[17242] = 8'h0e ;
            rom[17243] = 8'hfb ;
            rom[17244] = 8'h00 ;
            rom[17245] = 8'he6 ;
            rom[17246] = 8'he9 ;
            rom[17247] = 8'hf5 ;
            rom[17248] = 8'hf1 ;
            rom[17249] = 8'hf8 ;
            rom[17250] = 8'h04 ;
            rom[17251] = 8'h03 ;
            rom[17252] = 8'h11 ;
            rom[17253] = 8'h0e ;
            rom[17254] = 8'he5 ;
            rom[17255] = 8'hfe ;
            rom[17256] = 8'h17 ;
            rom[17257] = 8'h23 ;
            rom[17258] = 8'h20 ;
            rom[17259] = 8'hee ;
            rom[17260] = 8'h13 ;
            rom[17261] = 8'hfa ;
            rom[17262] = 8'hea ;
            rom[17263] = 8'hd2 ;
            rom[17264] = 8'h15 ;
            rom[17265] = 8'h01 ;
            rom[17266] = 8'hf5 ;
            rom[17267] = 8'h0f ;
            rom[17268] = 8'hf0 ;
            rom[17269] = 8'h0a ;
            rom[17270] = 8'hec ;
            rom[17271] = 8'he6 ;
            rom[17272] = 8'h04 ;
            rom[17273] = 8'he2 ;
            rom[17274] = 8'hfc ;
            rom[17275] = 8'hf9 ;
            rom[17276] = 8'hf5 ;
            rom[17277] = 8'hfd ;
            rom[17278] = 8'hd2 ;
            rom[17279] = 8'hfc ;
            rom[17280] = 8'h11 ;
            rom[17281] = 8'hfd ;
            rom[17282] = 8'hf0 ;
            rom[17283] = 8'hfa ;
            rom[17284] = 8'he3 ;
            rom[17285] = 8'hdc ;
            rom[17286] = 8'h03 ;
            rom[17287] = 8'he5 ;
            rom[17288] = 8'h13 ;
            rom[17289] = 8'hd7 ;
            rom[17290] = 8'h24 ;
            rom[17291] = 8'h33 ;
            rom[17292] = 8'hec ;
            rom[17293] = 8'h09 ;
            rom[17294] = 8'h17 ;
            rom[17295] = 8'hf2 ;
            rom[17296] = 8'he3 ;
            rom[17297] = 8'h06 ;
            rom[17298] = 8'hee ;
            rom[17299] = 8'h0d ;
            rom[17300] = 8'h07 ;
            rom[17301] = 8'h08 ;
            rom[17302] = 8'hc4 ;
            rom[17303] = 8'hbf ;
            rom[17304] = 8'hf9 ;
            rom[17305] = 8'h08 ;
            rom[17306] = 8'hfd ;
            rom[17307] = 8'hd2 ;
            rom[17308] = 8'h26 ;
            rom[17309] = 8'h00 ;
            rom[17310] = 8'h05 ;
            rom[17311] = 8'hef ;
            rom[17312] = 8'h14 ;
            rom[17313] = 8'h05 ;
            rom[17314] = 8'h0d ;
            rom[17315] = 8'hfd ;
            rom[17316] = 8'hfc ;
            rom[17317] = 8'h01 ;
            rom[17318] = 8'hda ;
            rom[17319] = 8'hee ;
            rom[17320] = 8'hfe ;
            rom[17321] = 8'h06 ;
            rom[17322] = 8'h14 ;
            rom[17323] = 8'hef ;
            rom[17324] = 8'h05 ;
            rom[17325] = 8'hfe ;
            rom[17326] = 8'h07 ;
            rom[17327] = 8'h04 ;
            rom[17328] = 8'heb ;
            rom[17329] = 8'h19 ;
            rom[17330] = 8'hd8 ;
            rom[17331] = 8'hd4 ;
            rom[17332] = 8'hfb ;
            rom[17333] = 8'h18 ;
            rom[17334] = 8'hfe ;
            rom[17335] = 8'hec ;
            rom[17336] = 8'h02 ;
            rom[17337] = 8'h00 ;
            rom[17338] = 8'h02 ;
            rom[17339] = 8'hed ;
            rom[17340] = 8'h24 ;
            rom[17341] = 8'hfb ;
            rom[17342] = 8'hea ;
            rom[17343] = 8'hf6 ;
            rom[17344] = 8'h0f ;
            rom[17345] = 8'hf7 ;
            rom[17346] = 8'h0e ;
            rom[17347] = 8'h06 ;
            rom[17348] = 8'he8 ;
            rom[17349] = 8'hf8 ;
            rom[17350] = 8'h00 ;
            rom[17351] = 8'hec ;
            rom[17352] = 8'hff ;
            rom[17353] = 8'hf7 ;
            rom[17354] = 8'h0c ;
            rom[17355] = 8'h0b ;
            rom[17356] = 8'h03 ;
            rom[17357] = 8'hff ;
            rom[17358] = 8'h0c ;
            rom[17359] = 8'he2 ;
            rom[17360] = 8'h06 ;
            rom[17361] = 8'hc3 ;
            rom[17362] = 8'he4 ;
            rom[17363] = 8'hf5 ;
            rom[17364] = 8'h07 ;
            rom[17365] = 8'h25 ;
            rom[17366] = 8'he4 ;
            rom[17367] = 8'hfe ;
            rom[17368] = 8'h0a ;
            rom[17369] = 8'h0d ;
            rom[17370] = 8'hed ;
            rom[17371] = 8'h05 ;
            rom[17372] = 8'h0f ;
            rom[17373] = 8'h1c ;
            rom[17374] = 8'h02 ;
            rom[17375] = 8'hdc ;
            rom[17376] = 8'h0c ;
            rom[17377] = 8'h0a ;
            rom[17378] = 8'h01 ;
            rom[17379] = 8'h02 ;
            rom[17380] = 8'hf9 ;
            rom[17381] = 8'h18 ;
            rom[17382] = 8'hdb ;
            rom[17383] = 8'hf1 ;
            rom[17384] = 8'h2d ;
            rom[17385] = 8'h07 ;
            rom[17386] = 8'hf6 ;
            rom[17387] = 8'h05 ;
            rom[17388] = 8'hed ;
            rom[17389] = 8'he6 ;
            rom[17390] = 8'hf1 ;
            rom[17391] = 8'h10 ;
            rom[17392] = 8'hc8 ;
            rom[17393] = 8'hf7 ;
            rom[17394] = 8'hec ;
            rom[17395] = 8'he5 ;
            rom[17396] = 8'he8 ;
            rom[17397] = 8'h4a ;
            rom[17398] = 8'h03 ;
            rom[17399] = 8'hfe ;
            rom[17400] = 8'h06 ;
            rom[17401] = 8'h0f ;
            rom[17402] = 8'hf6 ;
            rom[17403] = 8'he6 ;
            rom[17404] = 8'hd6 ;
            rom[17405] = 8'hfe ;
            rom[17406] = 8'h20 ;
            rom[17407] = 8'hf1 ;
            rom[17408] = 8'h02 ;
            rom[17409] = 8'h0a ;
            rom[17410] = 8'h07 ;
            rom[17411] = 8'hff ;
            rom[17412] = 8'hf4 ;
            rom[17413] = 8'hed ;
            rom[17414] = 8'h05 ;
            rom[17415] = 8'h20 ;
            rom[17416] = 8'h11 ;
            rom[17417] = 8'h13 ;
            rom[17418] = 8'hee ;
            rom[17419] = 8'hf1 ;
            rom[17420] = 8'hf5 ;
            rom[17421] = 8'h07 ;
            rom[17422] = 8'hdc ;
            rom[17423] = 8'hfe ;
            rom[17424] = 8'h09 ;
            rom[17425] = 8'hec ;
            rom[17426] = 8'hfa ;
            rom[17427] = 8'h05 ;
            rom[17428] = 8'h0c ;
            rom[17429] = 8'h05 ;
            rom[17430] = 8'hde ;
            rom[17431] = 8'hf1 ;
            rom[17432] = 8'hf1 ;
            rom[17433] = 8'hfb ;
            rom[17434] = 8'he9 ;
            rom[17435] = 8'h16 ;
            rom[17436] = 8'he5 ;
            rom[17437] = 8'h0d ;
            rom[17438] = 8'h0c ;
            rom[17439] = 8'h08 ;
            rom[17440] = 8'h08 ;
            rom[17441] = 8'h21 ;
            rom[17442] = 8'h01 ;
            rom[17443] = 8'h0c ;
            rom[17444] = 8'h0b ;
            rom[17445] = 8'hdf ;
            rom[17446] = 8'hd9 ;
            rom[17447] = 8'hf8 ;
            rom[17448] = 8'h18 ;
            rom[17449] = 8'hfc ;
            rom[17450] = 8'h09 ;
            rom[17451] = 8'hf2 ;
            rom[17452] = 8'hea ;
            rom[17453] = 8'hf9 ;
            rom[17454] = 8'hf3 ;
            rom[17455] = 8'h14 ;
            rom[17456] = 8'he5 ;
            rom[17457] = 8'he9 ;
            rom[17458] = 8'hf0 ;
            rom[17459] = 8'hcb ;
            rom[17460] = 8'h13 ;
            rom[17461] = 8'h10 ;
            rom[17462] = 8'hf0 ;
            rom[17463] = 8'hee ;
            rom[17464] = 8'h12 ;
            rom[17465] = 8'h12 ;
            rom[17466] = 8'h03 ;
            rom[17467] = 8'hed ;
            rom[17468] = 8'hf7 ;
            rom[17469] = 8'hf3 ;
            rom[17470] = 8'h0a ;
            rom[17471] = 8'h0a ;
            rom[17472] = 8'hf9 ;
            rom[17473] = 8'h08 ;
            rom[17474] = 8'hfb ;
            rom[17475] = 8'h07 ;
            rom[17476] = 8'h04 ;
            rom[17477] = 8'h04 ;
            rom[17478] = 8'h17 ;
            rom[17479] = 8'h1f ;
            rom[17480] = 8'hf8 ;
            rom[17481] = 8'h2f ;
            rom[17482] = 8'hef ;
            rom[17483] = 8'hf4 ;
            rom[17484] = 8'h08 ;
            rom[17485] = 8'h00 ;
            rom[17486] = 8'h1d ;
            rom[17487] = 8'h1f ;
            rom[17488] = 8'hec ;
            rom[17489] = 8'hf8 ;
            rom[17490] = 8'h0b ;
            rom[17491] = 8'h11 ;
            rom[17492] = 8'hf5 ;
            rom[17493] = 8'he9 ;
            rom[17494] = 8'he1 ;
            rom[17495] = 8'hee ;
            rom[17496] = 8'he3 ;
            rom[17497] = 8'hff ;
            rom[17498] = 8'h01 ;
            rom[17499] = 8'hd1 ;
            rom[17500] = 8'h10 ;
            rom[17501] = 8'he6 ;
            rom[17502] = 8'he2 ;
            rom[17503] = 8'he8 ;
            rom[17504] = 8'h13 ;
            rom[17505] = 8'he9 ;
            rom[17506] = 8'hf6 ;
            rom[17507] = 8'h02 ;
            rom[17508] = 8'hfc ;
            rom[17509] = 8'hf8 ;
            rom[17510] = 8'h08 ;
            rom[17511] = 8'hef ;
            rom[17512] = 8'hdd ;
            rom[17513] = 8'h1f ;
            rom[17514] = 8'h00 ;
            rom[17515] = 8'hf4 ;
            rom[17516] = 8'hf1 ;
            rom[17517] = 8'h06 ;
            rom[17518] = 8'hea ;
            rom[17519] = 8'hfe ;
            rom[17520] = 8'hfb ;
            rom[17521] = 8'h09 ;
            rom[17522] = 8'hec ;
            rom[17523] = 8'h10 ;
            rom[17524] = 8'h01 ;
            rom[17525] = 8'hf2 ;
            rom[17526] = 8'h08 ;
            rom[17527] = 8'h05 ;
            rom[17528] = 8'h07 ;
            rom[17529] = 8'hd3 ;
            rom[17530] = 8'h1a ;
            rom[17531] = 8'hf7 ;
            rom[17532] = 8'h22 ;
            rom[17533] = 8'hf4 ;
            rom[17534] = 8'hf1 ;
            rom[17535] = 8'h18 ;
            rom[17536] = 8'hef ;
            rom[17537] = 8'h07 ;
            rom[17538] = 8'h01 ;
            rom[17539] = 8'h14 ;
            rom[17540] = 8'h08 ;
            rom[17541] = 8'he5 ;
            rom[17542] = 8'h1a ;
            rom[17543] = 8'h0d ;
            rom[17544] = 8'h05 ;
            rom[17545] = 8'h06 ;
            rom[17546] = 8'h1c ;
            rom[17547] = 8'h02 ;
            rom[17548] = 8'he0 ;
            rom[17549] = 8'he2 ;
            rom[17550] = 8'hfe ;
            rom[17551] = 8'h05 ;
            rom[17552] = 8'hfb ;
            rom[17553] = 8'hfc ;
            rom[17554] = 8'h11 ;
            rom[17555] = 8'h22 ;
            rom[17556] = 8'hed ;
            rom[17557] = 8'h0f ;
            rom[17558] = 8'he2 ;
            rom[17559] = 8'h32 ;
            rom[17560] = 8'h02 ;
            rom[17561] = 8'h00 ;
            rom[17562] = 8'h13 ;
            rom[17563] = 8'hf2 ;
            rom[17564] = 8'hc3 ;
            rom[17565] = 8'h15 ;
            rom[17566] = 8'h0c ;
            rom[17567] = 8'he7 ;
            rom[17568] = 8'h10 ;
            rom[17569] = 8'hf0 ;
            rom[17570] = 8'h01 ;
            rom[17571] = 8'he6 ;
            rom[17572] = 8'hfb ;
            rom[17573] = 8'hf7 ;
            rom[17574] = 8'he4 ;
            rom[17575] = 8'h01 ;
            rom[17576] = 8'h18 ;
            rom[17577] = 8'h18 ;
            rom[17578] = 8'h12 ;
            rom[17579] = 8'h01 ;
            rom[17580] = 8'hd8 ;
            rom[17581] = 8'he3 ;
            rom[17582] = 8'h05 ;
            rom[17583] = 8'hd0 ;
            rom[17584] = 8'h00 ;
            rom[17585] = 8'h0a ;
            rom[17586] = 8'he5 ;
            rom[17587] = 8'hd8 ;
            rom[17588] = 8'hf7 ;
            rom[17589] = 8'h12 ;
            rom[17590] = 8'hfe ;
            rom[17591] = 8'hdc ;
            rom[17592] = 8'hf9 ;
            rom[17593] = 8'h09 ;
            rom[17594] = 8'h08 ;
            rom[17595] = 8'hf4 ;
            rom[17596] = 8'hec ;
            rom[17597] = 8'h08 ;
            rom[17598] = 8'hee ;
            rom[17599] = 8'hf5 ;
            rom[17600] = 8'hfa ;
            rom[17601] = 8'h1a ;
            rom[17602] = 8'h05 ;
            rom[17603] = 8'h09 ;
            rom[17604] = 8'hcd ;
            rom[17605] = 8'hf7 ;
            rom[17606] = 8'hfc ;
            rom[17607] = 8'he9 ;
            rom[17608] = 8'hc2 ;
            rom[17609] = 8'h04 ;
            rom[17610] = 8'heb ;
            rom[17611] = 8'h10 ;
            rom[17612] = 8'h18 ;
            rom[17613] = 8'h11 ;
            rom[17614] = 8'h05 ;
            rom[17615] = 8'h0e ;
            rom[17616] = 8'h9f ;
            rom[17617] = 8'heb ;
            rom[17618] = 8'h24 ;
            rom[17619] = 8'hf4 ;
            rom[17620] = 8'hd8 ;
            rom[17621] = 8'h28 ;
            rom[17622] = 8'h03 ;
            rom[17623] = 8'he4 ;
            rom[17624] = 8'hfa ;
            rom[17625] = 8'he8 ;
            rom[17626] = 8'h14 ;
            rom[17627] = 8'h09 ;
            rom[17628] = 8'h03 ;
            rom[17629] = 8'hd5 ;
            rom[17630] = 8'hf0 ;
            rom[17631] = 8'hf3 ;
            rom[17632] = 8'h11 ;
            rom[17633] = 8'hd0 ;
            rom[17634] = 8'h16 ;
            rom[17635] = 8'hd1 ;
            rom[17636] = 8'hff ;
            rom[17637] = 8'h10 ;
            rom[17638] = 8'h00 ;
            rom[17639] = 8'hfa ;
            rom[17640] = 8'hf6 ;
            rom[17641] = 8'h08 ;
            rom[17642] = 8'hce ;
            rom[17643] = 8'h1a ;
            rom[17644] = 8'hef ;
            rom[17645] = 8'h03 ;
            rom[17646] = 8'hdf ;
            rom[17647] = 8'hf3 ;
            rom[17648] = 8'h0f ;
            rom[17649] = 8'hea ;
            rom[17650] = 8'hfa ;
            rom[17651] = 8'h01 ;
            rom[17652] = 8'hfd ;
            rom[17653] = 8'h00 ;
            rom[17654] = 8'hfc ;
            rom[17655] = 8'hf3 ;
            rom[17656] = 8'h30 ;
            rom[17657] = 8'h2a ;
            rom[17658] = 8'hf6 ;
            rom[17659] = 8'hfa ;
            rom[17660] = 8'h00 ;
            rom[17661] = 8'h11 ;
            rom[17662] = 8'h13 ;
            rom[17663] = 8'hf2 ;
            rom[17664] = 8'h18 ;
            rom[17665] = 8'h0b ;
            rom[17666] = 8'h04 ;
            rom[17667] = 8'h19 ;
            rom[17668] = 8'hf9 ;
            rom[17669] = 8'hfb ;
            rom[17670] = 8'h05 ;
            rom[17671] = 8'hfe ;
            rom[17672] = 8'h02 ;
            rom[17673] = 8'h1a ;
            rom[17674] = 8'heb ;
            rom[17675] = 8'h02 ;
            rom[17676] = 8'h1c ;
            rom[17677] = 8'h0a ;
            rom[17678] = 8'hcc ;
            rom[17679] = 8'hed ;
            rom[17680] = 8'he0 ;
            rom[17681] = 8'h14 ;
            rom[17682] = 8'h1b ;
            rom[17683] = 8'h17 ;
            rom[17684] = 8'hfa ;
            rom[17685] = 8'hd2 ;
            rom[17686] = 8'hf3 ;
            rom[17687] = 8'h15 ;
            rom[17688] = 8'hf7 ;
            rom[17689] = 8'hf2 ;
            rom[17690] = 8'h14 ;
            rom[17691] = 8'h0c ;
            rom[17692] = 8'h08 ;
            rom[17693] = 8'he4 ;
            rom[17694] = 8'h0d ;
            rom[17695] = 8'h12 ;
            rom[17696] = 8'he8 ;
            rom[17697] = 8'h12 ;
            rom[17698] = 8'h19 ;
            rom[17699] = 8'hfa ;
            rom[17700] = 8'h19 ;
            rom[17701] = 8'hee ;
            rom[17702] = 8'hdb ;
            rom[17703] = 8'h03 ;
            rom[17704] = 8'h1b ;
            rom[17705] = 8'h26 ;
            rom[17706] = 8'h17 ;
            rom[17707] = 8'hf3 ;
            rom[17708] = 8'h02 ;
            rom[17709] = 8'h08 ;
            rom[17710] = 8'h0d ;
            rom[17711] = 8'h02 ;
            rom[17712] = 8'he8 ;
            rom[17713] = 8'h0f ;
            rom[17714] = 8'hc5 ;
            rom[17715] = 8'h0f ;
            rom[17716] = 8'he6 ;
            rom[17717] = 8'he5 ;
            rom[17718] = 8'hfe ;
            rom[17719] = 8'he6 ;
            rom[17720] = 8'h0a ;
            rom[17721] = 8'hfc ;
            rom[17722] = 8'hfc ;
            rom[17723] = 8'hf8 ;
            rom[17724] = 8'h21 ;
            rom[17725] = 8'h0a ;
            rom[17726] = 8'hf0 ;
            rom[17727] = 8'h0c ;
            rom[17728] = 8'hfe ;
            rom[17729] = 8'hd5 ;
            rom[17730] = 8'h15 ;
            rom[17731] = 8'hfa ;
            rom[17732] = 8'hf9 ;
            rom[17733] = 8'he9 ;
            rom[17734] = 8'hed ;
            rom[17735] = 8'hf2 ;
            rom[17736] = 8'h0d ;
            rom[17737] = 8'h02 ;
            rom[17738] = 8'h17 ;
            rom[17739] = 8'h30 ;
            rom[17740] = 8'h1a ;
            rom[17741] = 8'h0e ;
            rom[17742] = 8'h04 ;
            rom[17743] = 8'hf3 ;
            rom[17744] = 8'hf4 ;
            rom[17745] = 8'he1 ;
            rom[17746] = 8'hfd ;
            rom[17747] = 8'h06 ;
            rom[17748] = 8'he1 ;
            rom[17749] = 8'hf5 ;
            rom[17750] = 8'h00 ;
            rom[17751] = 8'hf2 ;
            rom[17752] = 8'h10 ;
            rom[17753] = 8'heb ;
            rom[17754] = 8'hf6 ;
            rom[17755] = 8'h17 ;
            rom[17756] = 8'hf6 ;
            rom[17757] = 8'hd7 ;
            rom[17758] = 8'he5 ;
            rom[17759] = 8'h00 ;
            rom[17760] = 8'he9 ;
            rom[17761] = 8'he0 ;
            rom[17762] = 8'hfc ;
            rom[17763] = 8'hf2 ;
            rom[17764] = 8'h21 ;
            rom[17765] = 8'heb ;
            rom[17766] = 8'hfb ;
            rom[17767] = 8'he8 ;
            rom[17768] = 8'hfa ;
            rom[17769] = 8'he8 ;
            rom[17770] = 8'he7 ;
            rom[17771] = 8'h08 ;
            rom[17772] = 8'h00 ;
            rom[17773] = 8'hfd ;
            rom[17774] = 8'h0a ;
            rom[17775] = 8'h08 ;
            rom[17776] = 8'hca ;
            rom[17777] = 8'hea ;
            rom[17778] = 8'h05 ;
            rom[17779] = 8'hff ;
            rom[17780] = 8'hfe ;
            rom[17781] = 8'h11 ;
            rom[17782] = 8'he1 ;
            rom[17783] = 8'hfd ;
            rom[17784] = 8'h14 ;
            rom[17785] = 8'heb ;
            rom[17786] = 8'h13 ;
            rom[17787] = 8'hee ;
            rom[17788] = 8'h12 ;
            rom[17789] = 8'h14 ;
            rom[17790] = 8'h18 ;
            rom[17791] = 8'h03 ;
            rom[17792] = 8'h05 ;
            rom[17793] = 8'hce ;
            rom[17794] = 8'hf7 ;
            rom[17795] = 8'heb ;
            rom[17796] = 8'hfc ;
            rom[17797] = 8'h19 ;
            rom[17798] = 8'h13 ;
            rom[17799] = 8'hee ;
            rom[17800] = 8'h0f ;
            rom[17801] = 8'h1d ;
            rom[17802] = 8'h16 ;
            rom[17803] = 8'h27 ;
            rom[17804] = 8'hf8 ;
            rom[17805] = 8'h01 ;
            rom[17806] = 8'hda ;
            rom[17807] = 8'hf1 ;
            rom[17808] = 8'h0d ;
            rom[17809] = 8'hf6 ;
            rom[17810] = 8'hdb ;
            rom[17811] = 8'hde ;
            rom[17812] = 8'h07 ;
            rom[17813] = 8'h0f ;
            rom[17814] = 8'h0b ;
            rom[17815] = 8'h1a ;
            rom[17816] = 8'hfa ;
            rom[17817] = 8'he1 ;
            rom[17818] = 8'h1b ;
            rom[17819] = 8'hde ;
            rom[17820] = 8'h20 ;
            rom[17821] = 8'hdd ;
            rom[17822] = 8'he8 ;
            rom[17823] = 8'h0d ;
            rom[17824] = 8'h00 ;
            rom[17825] = 8'h01 ;
            rom[17826] = 8'he0 ;
            rom[17827] = 8'heb ;
            rom[17828] = 8'h03 ;
            rom[17829] = 8'h03 ;
            rom[17830] = 8'h05 ;
            rom[17831] = 8'h1c ;
            rom[17832] = 8'hdb ;
            rom[17833] = 8'h09 ;
            rom[17834] = 8'hf5 ;
            rom[17835] = 8'hff ;
            rom[17836] = 8'he9 ;
            rom[17837] = 8'hf8 ;
            rom[17838] = 8'h25 ;
            rom[17839] = 8'hdf ;
            rom[17840] = 8'hf9 ;
            rom[17841] = 8'hd9 ;
            rom[17842] = 8'h03 ;
            rom[17843] = 8'hfa ;
            rom[17844] = 8'hf3 ;
            rom[17845] = 8'h04 ;
            rom[17846] = 8'hf8 ;
            rom[17847] = 8'h07 ;
            rom[17848] = 8'he6 ;
            rom[17849] = 8'h05 ;
            rom[17850] = 8'h15 ;
            rom[17851] = 8'hf8 ;
            rom[17852] = 8'hfc ;
            rom[17853] = 8'h14 ;
            rom[17854] = 8'h07 ;
            rom[17855] = 8'hea ;
            rom[17856] = 8'h00 ;
            rom[17857] = 8'hf8 ;
            rom[17858] = 8'h1e ;
            rom[17859] = 8'he7 ;
            rom[17860] = 8'hf6 ;
            rom[17861] = 8'h0b ;
            rom[17862] = 8'hd5 ;
            rom[17863] = 8'hfb ;
            rom[17864] = 8'hea ;
            rom[17865] = 8'hfd ;
            rom[17866] = 8'h2d ;
            rom[17867] = 8'h29 ;
            rom[17868] = 8'hee ;
            rom[17869] = 8'h1e ;
            rom[17870] = 8'h0f ;
            rom[17871] = 8'hf9 ;
            rom[17872] = 8'hd4 ;
            rom[17873] = 8'h08 ;
            rom[17874] = 8'h16 ;
            rom[17875] = 8'h0d ;
            rom[17876] = 8'he1 ;
            rom[17877] = 8'h05 ;
            rom[17878] = 8'hd8 ;
            rom[17879] = 8'hf4 ;
            rom[17880] = 8'h22 ;
            rom[17881] = 8'h1d ;
            rom[17882] = 8'hdf ;
            rom[17883] = 8'h04 ;
            rom[17884] = 8'h03 ;
            rom[17885] = 8'hcc ;
            rom[17886] = 8'he7 ;
            rom[17887] = 8'h19 ;
            rom[17888] = 8'hf8 ;
            rom[17889] = 8'hed ;
            rom[17890] = 8'hec ;
            rom[17891] = 8'hd4 ;
            rom[17892] = 8'h03 ;
            rom[17893] = 8'hfd ;
            rom[17894] = 8'h0f ;
            rom[17895] = 8'h0b ;
            rom[17896] = 8'hec ;
            rom[17897] = 8'h0c ;
            rom[17898] = 8'hfb ;
            rom[17899] = 8'h01 ;
            rom[17900] = 8'h12 ;
            rom[17901] = 8'he2 ;
            rom[17902] = 8'h14 ;
            rom[17903] = 8'hf9 ;
            rom[17904] = 8'hd9 ;
            rom[17905] = 8'h12 ;
            rom[17906] = 8'h19 ;
            rom[17907] = 8'h17 ;
            rom[17908] = 8'h0c ;
            rom[17909] = 8'h1c ;
            rom[17910] = 8'he4 ;
            rom[17911] = 8'hf8 ;
            rom[17912] = 8'h13 ;
            rom[17913] = 8'hf3 ;
            rom[17914] = 8'h0b ;
            rom[17915] = 8'h08 ;
            rom[17916] = 8'h15 ;
            rom[17917] = 8'h13 ;
            rom[17918] = 8'hfe ;
            rom[17919] = 8'he8 ;
            rom[17920] = 8'hf2 ;
            rom[17921] = 8'hd0 ;
            rom[17922] = 8'hf6 ;
            rom[17923] = 8'h0d ;
            rom[17924] = 8'hf5 ;
            rom[17925] = 8'hfd ;
            rom[17926] = 8'h1e ;
            rom[17927] = 8'h12 ;
            rom[17928] = 8'h05 ;
            rom[17929] = 8'h17 ;
            rom[17930] = 8'h06 ;
            rom[17931] = 8'h04 ;
            rom[17932] = 8'h1d ;
            rom[17933] = 8'h04 ;
            rom[17934] = 8'hea ;
            rom[17935] = 8'hf4 ;
            rom[17936] = 8'h01 ;
            rom[17937] = 8'h07 ;
            rom[17938] = 8'h21 ;
            rom[17939] = 8'h24 ;
            rom[17940] = 8'he8 ;
            rom[17941] = 8'h1f ;
            rom[17942] = 8'he9 ;
            rom[17943] = 8'h13 ;
            rom[17944] = 8'h0e ;
            rom[17945] = 8'h0f ;
            rom[17946] = 8'hfb ;
            rom[17947] = 8'hdd ;
            rom[17948] = 8'hee ;
            rom[17949] = 8'he4 ;
            rom[17950] = 8'he3 ;
            rom[17951] = 8'he9 ;
            rom[17952] = 8'hf5 ;
            rom[17953] = 8'hb8 ;
            rom[17954] = 8'hf0 ;
            rom[17955] = 8'h14 ;
            rom[17956] = 8'h0c ;
            rom[17957] = 8'hef ;
            rom[17958] = 8'h06 ;
            rom[17959] = 8'he3 ;
            rom[17960] = 8'hf5 ;
            rom[17961] = 8'h3b ;
            rom[17962] = 8'h1a ;
            rom[17963] = 8'hfd ;
            rom[17964] = 8'h05 ;
            rom[17965] = 8'h03 ;
            rom[17966] = 8'he4 ;
            rom[17967] = 8'h02 ;
            rom[17968] = 8'hed ;
            rom[17969] = 8'hf3 ;
            rom[17970] = 8'h13 ;
            rom[17971] = 8'heb ;
            rom[17972] = 8'h09 ;
            rom[17973] = 8'h20 ;
            rom[17974] = 8'h09 ;
            rom[17975] = 8'hd2 ;
            rom[17976] = 8'hec ;
            rom[17977] = 8'he2 ;
            rom[17978] = 8'h08 ;
            rom[17979] = 8'hec ;
            rom[17980] = 8'h07 ;
            rom[17981] = 8'h14 ;
            rom[17982] = 8'hf1 ;
            rom[17983] = 8'hfe ;
            rom[17984] = 8'hf9 ;
            rom[17985] = 8'hef ;
            rom[17986] = 8'h08 ;
            rom[17987] = 8'h2a ;
            rom[17988] = 8'hd4 ;
            rom[17989] = 8'h13 ;
            rom[17990] = 8'hfa ;
            rom[17991] = 8'hf6 ;
            rom[17992] = 8'hd6 ;
            rom[17993] = 8'h0d ;
            rom[17994] = 8'h0b ;
            rom[17995] = 8'h17 ;
            rom[17996] = 8'hfb ;
            rom[17997] = 8'h11 ;
            rom[17998] = 8'h12 ;
            rom[17999] = 8'h12 ;
            rom[18000] = 8'hb5 ;
            rom[18001] = 8'hf4 ;
            rom[18002] = 8'h0a ;
            rom[18003] = 8'hf8 ;
            rom[18004] = 8'he6 ;
            rom[18005] = 8'h17 ;
            rom[18006] = 8'hf7 ;
            rom[18007] = 8'hf3 ;
            rom[18008] = 8'hf1 ;
            rom[18009] = 8'he9 ;
            rom[18010] = 8'h17 ;
            rom[18011] = 8'hff ;
            rom[18012] = 8'h11 ;
            rom[18013] = 8'hd3 ;
            rom[18014] = 8'hee ;
            rom[18015] = 8'hf3 ;
            rom[18016] = 8'h0c ;
            rom[18017] = 8'hda ;
            rom[18018] = 8'h17 ;
            rom[18019] = 8'hdb ;
            rom[18020] = 8'h00 ;
            rom[18021] = 8'h11 ;
            rom[18022] = 8'hf8 ;
            rom[18023] = 8'h09 ;
            rom[18024] = 8'hfe ;
            rom[18025] = 8'h07 ;
            rom[18026] = 8'hd0 ;
            rom[18027] = 8'h10 ;
            rom[18028] = 8'hfe ;
            rom[18029] = 8'h06 ;
            rom[18030] = 8'hf4 ;
            rom[18031] = 8'h04 ;
            rom[18032] = 8'hfb ;
            rom[18033] = 8'hed ;
            rom[18034] = 8'hfc ;
            rom[18035] = 8'hf7 ;
            rom[18036] = 8'h10 ;
            rom[18037] = 8'h03 ;
            rom[18038] = 8'he3 ;
            rom[18039] = 8'hf6 ;
            rom[18040] = 8'h11 ;
            rom[18041] = 8'hfd ;
            rom[18042] = 8'h08 ;
            rom[18043] = 8'h02 ;
            rom[18044] = 8'h0c ;
            rom[18045] = 8'h07 ;
            rom[18046] = 8'h12 ;
            rom[18047] = 8'h0a ;
            rom[18048] = 8'h0e ;
            rom[18049] = 8'hd8 ;
            rom[18050] = 8'hfc ;
            rom[18051] = 8'hd2 ;
            rom[18052] = 8'hdd ;
            rom[18053] = 8'h04 ;
            rom[18054] = 8'hed ;
            rom[18055] = 8'h00 ;
            rom[18056] = 8'he5 ;
            rom[18057] = 8'h0b ;
            rom[18058] = 8'h09 ;
            rom[18059] = 8'h12 ;
            rom[18060] = 8'hf7 ;
            rom[18061] = 8'h03 ;
            rom[18062] = 8'h17 ;
            rom[18063] = 8'hfd ;
            rom[18064] = 8'he0 ;
            rom[18065] = 8'hd9 ;
            rom[18066] = 8'h05 ;
            rom[18067] = 8'he4 ;
            rom[18068] = 8'hd0 ;
            rom[18069] = 8'hff ;
            rom[18070] = 8'h06 ;
            rom[18071] = 8'h1a ;
            rom[18072] = 8'h08 ;
            rom[18073] = 8'hc1 ;
            rom[18074] = 8'h20 ;
            rom[18075] = 8'hf8 ;
            rom[18076] = 8'h19 ;
            rom[18077] = 8'hc1 ;
            rom[18078] = 8'he3 ;
            rom[18079] = 8'hf4 ;
            rom[18080] = 8'hfd ;
            rom[18081] = 8'hd2 ;
            rom[18082] = 8'h15 ;
            rom[18083] = 8'hda ;
            rom[18084] = 8'h04 ;
            rom[18085] = 8'hfc ;
            rom[18086] = 8'h10 ;
            rom[18087] = 8'hf8 ;
            rom[18088] = 8'h05 ;
            rom[18089] = 8'h25 ;
            rom[18090] = 8'hd6 ;
            rom[18091] = 8'h0d ;
            rom[18092] = 8'h12 ;
            rom[18093] = 8'h05 ;
            rom[18094] = 8'h12 ;
            rom[18095] = 8'he7 ;
            rom[18096] = 8'h14 ;
            rom[18097] = 8'he7 ;
            rom[18098] = 8'h19 ;
            rom[18099] = 8'h06 ;
            rom[18100] = 8'h12 ;
            rom[18101] = 8'hf5 ;
            rom[18102] = 8'hfa ;
            rom[18103] = 8'h08 ;
            rom[18104] = 8'h0e ;
            rom[18105] = 8'h01 ;
            rom[18106] = 8'h2c ;
            rom[18107] = 8'hec ;
            rom[18108] = 8'h16 ;
            rom[18109] = 8'hf0 ;
            rom[18110] = 8'h07 ;
            rom[18111] = 8'h0d ;
            rom[18112] = 8'h01 ;
            rom[18113] = 8'hf4 ;
            rom[18114] = 8'h00 ;
            rom[18115] = 8'hec ;
            rom[18116] = 8'hdc ;
            rom[18117] = 8'heb ;
            rom[18118] = 8'hf0 ;
            rom[18119] = 8'h04 ;
            rom[18120] = 8'hea ;
            rom[18121] = 8'h0b ;
            rom[18122] = 8'h24 ;
            rom[18123] = 8'h12 ;
            rom[18124] = 8'hf5 ;
            rom[18125] = 8'h0e ;
            rom[18126] = 8'h08 ;
            rom[18127] = 8'h15 ;
            rom[18128] = 8'hc4 ;
            rom[18129] = 8'hf5 ;
            rom[18130] = 8'h1c ;
            rom[18131] = 8'h06 ;
            rom[18132] = 8'h89 ;
            rom[18133] = 8'hff ;
            rom[18134] = 8'h0d ;
            rom[18135] = 8'hf8 ;
            rom[18136] = 8'h01 ;
            rom[18137] = 8'h08 ;
            rom[18138] = 8'h07 ;
            rom[18139] = 8'h07 ;
            rom[18140] = 8'hfb ;
            rom[18141] = 8'hce ;
            rom[18142] = 8'he8 ;
            rom[18143] = 8'hf4 ;
            rom[18144] = 8'hec ;
            rom[18145] = 8'hf4 ;
            rom[18146] = 8'h06 ;
            rom[18147] = 8'hc5 ;
            rom[18148] = 8'hfd ;
            rom[18149] = 8'hde ;
            rom[18150] = 8'h16 ;
            rom[18151] = 8'h0e ;
            rom[18152] = 8'hdb ;
            rom[18153] = 8'h0b ;
            rom[18154] = 8'he3 ;
            rom[18155] = 8'h09 ;
            rom[18156] = 8'hfb ;
            rom[18157] = 8'he8 ;
            rom[18158] = 8'h03 ;
            rom[18159] = 8'h12 ;
            rom[18160] = 8'h1f ;
            rom[18161] = 8'hfe ;
            rom[18162] = 8'h03 ;
            rom[18163] = 8'h10 ;
            rom[18164] = 8'h1e ;
            rom[18165] = 8'h02 ;
            rom[18166] = 8'he6 ;
            rom[18167] = 8'hfa ;
            rom[18168] = 8'h0c ;
            rom[18169] = 8'hf2 ;
            rom[18170] = 8'h08 ;
            rom[18171] = 8'hdb ;
            rom[18172] = 8'h11 ;
            rom[18173] = 8'h1e ;
            rom[18174] = 8'hec ;
            rom[18175] = 8'hbb ;
            rom[18176] = 8'h0b ;
            rom[18177] = 8'hf5 ;
            rom[18178] = 8'h14 ;
            rom[18179] = 8'hfa ;
            rom[18180] = 8'he1 ;
            rom[18181] = 8'hf2 ;
            rom[18182] = 8'he6 ;
            rom[18183] = 8'hfa ;
            rom[18184] = 8'hf7 ;
            rom[18185] = 8'h02 ;
            rom[18186] = 8'h0e ;
            rom[18187] = 8'h0e ;
            rom[18188] = 8'h07 ;
            rom[18189] = 8'h1f ;
            rom[18190] = 8'he6 ;
            rom[18191] = 8'hf1 ;
            rom[18192] = 8'hf3 ;
            rom[18193] = 8'h06 ;
            rom[18194] = 8'h0b ;
            rom[18195] = 8'hfc ;
            rom[18196] = 8'h11 ;
            rom[18197] = 8'hfa ;
            rom[18198] = 8'hd8 ;
            rom[18199] = 8'heb ;
            rom[18200] = 8'hf9 ;
            rom[18201] = 8'heb ;
            rom[18202] = 8'hfc ;
            rom[18203] = 8'h0f ;
            rom[18204] = 8'heb ;
            rom[18205] = 8'hfa ;
            rom[18206] = 8'hdd ;
            rom[18207] = 8'h0f ;
            rom[18208] = 8'hf3 ;
            rom[18209] = 8'hfd ;
            rom[18210] = 8'hf0 ;
            rom[18211] = 8'h10 ;
            rom[18212] = 8'h18 ;
            rom[18213] = 8'he3 ;
            rom[18214] = 8'he4 ;
            rom[18215] = 8'he7 ;
            rom[18216] = 8'hf5 ;
            rom[18217] = 8'heb ;
            rom[18218] = 8'he7 ;
            rom[18219] = 8'hf5 ;
            rom[18220] = 8'h01 ;
            rom[18221] = 8'he8 ;
            rom[18222] = 8'hfa ;
            rom[18223] = 8'h0c ;
            rom[18224] = 8'hf1 ;
            rom[18225] = 8'h19 ;
            rom[18226] = 8'h06 ;
            rom[18227] = 8'hfe ;
            rom[18228] = 8'h09 ;
            rom[18229] = 8'h01 ;
            rom[18230] = 8'hf6 ;
            rom[18231] = 8'hd9 ;
            rom[18232] = 8'h11 ;
            rom[18233] = 8'hed ;
            rom[18234] = 8'h15 ;
            rom[18235] = 8'he3 ;
            rom[18236] = 8'h0b ;
            rom[18237] = 8'h0b ;
            rom[18238] = 8'h12 ;
            rom[18239] = 8'h08 ;
            rom[18240] = 8'h1b ;
            rom[18241] = 8'hef ;
            rom[18242] = 8'h0d ;
            rom[18243] = 8'he1 ;
            rom[18244] = 8'hec ;
            rom[18245] = 8'hee ;
            rom[18246] = 8'h19 ;
            rom[18247] = 8'he3 ;
            rom[18248] = 8'hfb ;
            rom[18249] = 8'h0f ;
            rom[18250] = 8'h0e ;
            rom[18251] = 8'hf6 ;
            rom[18252] = 8'h17 ;
            rom[18253] = 8'h24 ;
            rom[18254] = 8'h14 ;
            rom[18255] = 8'hc5 ;
            rom[18256] = 8'hee ;
            rom[18257] = 8'he7 ;
            rom[18258] = 8'hee ;
            rom[18259] = 8'h0c ;
            rom[18260] = 8'hf8 ;
            rom[18261] = 8'he5 ;
            rom[18262] = 8'hf5 ;
            rom[18263] = 8'hf9 ;
            rom[18264] = 8'h01 ;
            rom[18265] = 8'hef ;
            rom[18266] = 8'hf3 ;
            rom[18267] = 8'h08 ;
            rom[18268] = 8'hfb ;
            rom[18269] = 8'hd0 ;
            rom[18270] = 8'hfa ;
            rom[18271] = 8'h28 ;
            rom[18272] = 8'h0c ;
            rom[18273] = 8'hf0 ;
            rom[18274] = 8'h10 ;
            rom[18275] = 8'h0c ;
            rom[18276] = 8'h01 ;
            rom[18277] = 8'h38 ;
            rom[18278] = 8'hf2 ;
            rom[18279] = 8'hcc ;
            rom[18280] = 8'heb ;
            rom[18281] = 8'h14 ;
            rom[18282] = 8'hfd ;
            rom[18283] = 8'h00 ;
            rom[18284] = 8'h11 ;
            rom[18285] = 8'h00 ;
            rom[18286] = 8'hf9 ;
            rom[18287] = 8'he7 ;
            rom[18288] = 8'he4 ;
            rom[18289] = 8'hdd ;
            rom[18290] = 8'hc3 ;
            rom[18291] = 8'h0e ;
            rom[18292] = 8'h09 ;
            rom[18293] = 8'he8 ;
            rom[18294] = 8'h1c ;
            rom[18295] = 8'h10 ;
            rom[18296] = 8'h09 ;
            rom[18297] = 8'hea ;
            rom[18298] = 8'hf6 ;
            rom[18299] = 8'h0b ;
            rom[18300] = 8'hfb ;
            rom[18301] = 8'hed ;
            rom[18302] = 8'h04 ;
            rom[18303] = 8'h1b ;
            rom[18304] = 8'hf6 ;
            rom[18305] = 8'hf6 ;
            rom[18306] = 8'hf9 ;
            rom[18307] = 8'hdf ;
            rom[18308] = 8'hfd ;
            rom[18309] = 8'h06 ;
            rom[18310] = 8'h05 ;
            rom[18311] = 8'heb ;
            rom[18312] = 8'h0d ;
            rom[18313] = 8'hf8 ;
            rom[18314] = 8'h08 ;
            rom[18315] = 8'h11 ;
            rom[18316] = 8'hd9 ;
            rom[18317] = 8'hc6 ;
            rom[18318] = 8'hf9 ;
            rom[18319] = 8'he1 ;
            rom[18320] = 8'h0a ;
            rom[18321] = 8'he7 ;
            rom[18322] = 8'heb ;
            rom[18323] = 8'h01 ;
            rom[18324] = 8'h12 ;
            rom[18325] = 8'h2c ;
            rom[18326] = 8'h17 ;
            rom[18327] = 8'hf8 ;
            rom[18328] = 8'hf4 ;
            rom[18329] = 8'h0a ;
            rom[18330] = 8'h1e ;
            rom[18331] = 8'h07 ;
            rom[18332] = 8'h10 ;
            rom[18333] = 8'hef ;
            rom[18334] = 8'hd8 ;
            rom[18335] = 8'hfd ;
            rom[18336] = 8'hf5 ;
            rom[18337] = 8'hf4 ;
            rom[18338] = 8'hf2 ;
            rom[18339] = 8'hff ;
            rom[18340] = 8'h01 ;
            rom[18341] = 8'h21 ;
            rom[18342] = 8'hed ;
            rom[18343] = 8'h0a ;
            rom[18344] = 8'h16 ;
            rom[18345] = 8'hf9 ;
            rom[18346] = 8'h1b ;
            rom[18347] = 8'hf3 ;
            rom[18348] = 8'hfb ;
            rom[18349] = 8'h1b ;
            rom[18350] = 8'hff ;
            rom[18351] = 8'hfe ;
            rom[18352] = 8'he4 ;
            rom[18353] = 8'hea ;
            rom[18354] = 8'hfa ;
            rom[18355] = 8'hcd ;
            rom[18356] = 8'he8 ;
            rom[18357] = 8'h14 ;
            rom[18358] = 8'h02 ;
            rom[18359] = 8'h03 ;
            rom[18360] = 8'hee ;
            rom[18361] = 8'h1d ;
            rom[18362] = 8'hf5 ;
            rom[18363] = 8'hf5 ;
            rom[18364] = 8'hf4 ;
            rom[18365] = 8'h11 ;
            rom[18366] = 8'h08 ;
            rom[18367] = 8'hdc ;
            rom[18368] = 8'h0e ;
            rom[18369] = 8'hf4 ;
            rom[18370] = 8'hfd ;
            rom[18371] = 8'h11 ;
            rom[18372] = 8'he8 ;
            rom[18373] = 8'hf8 ;
            rom[18374] = 8'hfa ;
            rom[18375] = 8'h14 ;
            rom[18376] = 8'hfa ;
            rom[18377] = 8'hf7 ;
            rom[18378] = 8'h13 ;
            rom[18379] = 8'h0d ;
            rom[18380] = 8'h21 ;
            rom[18381] = 8'h07 ;
            rom[18382] = 8'h18 ;
            rom[18383] = 8'hd9 ;
            rom[18384] = 8'h05 ;
            rom[18385] = 8'hef ;
            rom[18386] = 8'h1e ;
            rom[18387] = 8'hf5 ;
            rom[18388] = 8'heb ;
            rom[18389] = 8'hfa ;
            rom[18390] = 8'hd3 ;
            rom[18391] = 8'h14 ;
            rom[18392] = 8'h19 ;
            rom[18393] = 8'h1e ;
            rom[18394] = 8'he3 ;
            rom[18395] = 8'h0a ;
            rom[18396] = 8'h17 ;
            rom[18397] = 8'he5 ;
            rom[18398] = 8'h18 ;
            rom[18399] = 8'hf4 ;
            rom[18400] = 8'h08 ;
            rom[18401] = 8'hf6 ;
            rom[18402] = 8'hf5 ;
            rom[18403] = 8'h07 ;
            rom[18404] = 8'h17 ;
            rom[18405] = 8'h1f ;
            rom[18406] = 8'h13 ;
            rom[18407] = 8'hd5 ;
            rom[18408] = 8'hf8 ;
            rom[18409] = 8'hef ;
            rom[18410] = 8'h0c ;
            rom[18411] = 8'h18 ;
            rom[18412] = 8'h1a ;
            rom[18413] = 8'h01 ;
            rom[18414] = 8'h0b ;
            rom[18415] = 8'hee ;
            rom[18416] = 8'he1 ;
            rom[18417] = 8'hdb ;
            rom[18418] = 8'he2 ;
            rom[18419] = 8'h18 ;
            rom[18420] = 8'h25 ;
            rom[18421] = 8'h10 ;
            rom[18422] = 8'h10 ;
            rom[18423] = 8'hfd ;
            rom[18424] = 8'h15 ;
            rom[18425] = 8'hf5 ;
            rom[18426] = 8'h03 ;
            rom[18427] = 8'hfb ;
            rom[18428] = 8'h19 ;
            rom[18429] = 8'hef ;
            rom[18430] = 8'h10 ;
            rom[18431] = 8'hfc ;
        end
    always
        @(*)
        begin
            data = rom[addr] ;
        end
endmodule



