
module weights_rom_dense_layer_2x_128_to_9 (
    input wire [10:0] addr, 
    output reg signed [7:0] data) ;
    reg signed [7:0] rom [0:1151] ; 
    initial
        begin
            rom[0] = 8'hce ;
            rom[1] = 8'hd2 ;
            rom[2] = 8'h29 ;
            rom[3] = 8'he6 ;
            rom[4] = 8'h37 ;
            rom[5] = 8'h35 ;
            rom[6] = 8'h40 ;
            rom[7] = 8'h38 ;
            rom[8] = 8'hc6 ;
            rom[9] = 8'hbc ;
            rom[10] = 8'h37 ;
            rom[11] = 8'h97 ;
            rom[12] = 8'h30 ;
            rom[13] = 8'h3e ;
            rom[14] = 8'h35 ;
            rom[15] = 8'h46 ;
            rom[16] = 8'h49 ;
            rom[17] = 8'hed ;
            rom[18] = 8'h95 ;
            rom[19] = 8'ha8 ;
            rom[20] = 8'h20 ;
            rom[21] = 8'had ;
            rom[22] = 8'hea ;
            rom[23] = 8'he0 ;
            rom[24] = 8'hcf ;
            rom[25] = 8'he5 ;
            rom[26] = 8'h2c ;
            rom[27] = 8'h15 ;
            rom[28] = 8'hd4 ;
            rom[29] = 8'h14 ;
            rom[30] = 8'hb2 ;
            rom[31] = 8'h35 ;
            rom[32] = 8'h15 ;
            rom[33] = 8'hd0 ;
            rom[34] = 8'h29 ;
            rom[35] = 8'hc6 ;
            rom[36] = 8'hf7 ;
            rom[37] = 8'h12 ;
            rom[38] = 8'hd6 ;
            rom[39] = 8'h30 ;
            rom[40] = 8'h41 ;
            rom[41] = 8'hfe ;
            rom[42] = 8'h40 ;
            rom[43] = 8'he3 ;
            rom[44] = 8'h05 ;
            rom[45] = 8'he1 ;
            rom[46] = 8'hf7 ;
            rom[47] = 8'h09 ;
            rom[48] = 8'h47 ;
            rom[49] = 8'hf2 ;
            rom[50] = 8'h31 ;
            rom[51] = 8'h03 ;
            rom[52] = 8'h2e ;
            rom[53] = 8'h43 ;
            rom[54] = 8'h3d ;
            rom[55] = 8'h35 ;
            rom[56] = 8'hd9 ;
            rom[57] = 8'hf4 ;
            rom[58] = 8'hcf ;
            rom[59] = 8'hed ;
            rom[60] = 8'hdf ;
            rom[61] = 8'h36 ;
            rom[62] = 8'hea ;
            rom[63] = 8'he3 ;
            rom[64] = 8'hdc ;
            rom[65] = 8'he4 ;
            rom[66] = 8'h4c ;
            rom[67] = 8'hdb ;
            rom[68] = 8'h52 ;
            rom[69] = 8'heb ;
            rom[70] = 8'hde ;
            rom[71] = 8'h68 ;
            rom[72] = 8'hdf ;
            rom[73] = 8'hdd ;
            rom[74] = 8'hee ;
            rom[75] = 8'hf1 ;
            rom[76] = 8'he8 ;
            rom[77] = 8'he0 ;
            rom[78] = 8'hec ;
            rom[79] = 8'h56 ;
            rom[80] = 8'h00 ;
            rom[81] = 8'h05 ;
            rom[82] = 8'he7 ;
            rom[83] = 8'hea ;
            rom[84] = 8'hda ;
            rom[85] = 8'h2f ;
            rom[86] = 8'h40 ;
            rom[87] = 8'hc8 ;
            rom[88] = 8'he1 ;
            rom[89] = 8'h1f ;
            rom[90] = 8'hc3 ;
            rom[91] = 8'hb7 ;
            rom[92] = 8'h1c ;
            rom[93] = 8'h1e ;
            rom[94] = 8'h35 ;
            rom[95] = 8'h48 ;
            rom[96] = 8'hd8 ;
            rom[97] = 8'h36 ;
            rom[98] = 8'hcf ;
            rom[99] = 8'hca ;
            rom[100] = 8'he5 ;
            rom[101] = 8'h37 ;
            rom[102] = 8'he1 ;
            rom[103] = 8'h47 ;
            rom[104] = 8'hec ;
            rom[105] = 8'h3d ;
            rom[106] = 8'he0 ;
            rom[107] = 8'hef ;
            rom[108] = 8'h51 ;
            rom[109] = 8'h42 ;
            rom[110] = 8'h13 ;
            rom[111] = 8'h54 ;
            rom[112] = 8'h33 ;
            rom[113] = 8'hdd ;
            rom[114] = 8'h13 ;
            rom[115] = 8'hd4 ;
            rom[116] = 8'hd8 ;
            rom[117] = 8'hda ;
            rom[118] = 8'hd9 ;
            rom[119] = 8'hf0 ;
            rom[120] = 8'hc5 ;
            rom[121] = 8'hb6 ;
            rom[122] = 8'h30 ;
            rom[123] = 8'h31 ;
            rom[124] = 8'h3f ;
            rom[125] = 8'h32 ;
            rom[126] = 8'hb4 ;
            rom[127] = 8'h33 ;
            rom[128] = 8'hc9 ;
            rom[129] = 8'hd1 ;
            rom[130] = 8'haf ;
            rom[131] = 8'ha4 ;
            rom[132] = 8'h08 ;
            rom[133] = 8'hd3 ;
            rom[134] = 8'h1a ;
            rom[135] = 8'h17 ;
            rom[136] = 8'hd0 ;
            rom[137] = 8'h17 ;
            rom[138] = 8'hbd ;
            rom[139] = 8'h97 ;
            rom[140] = 8'hf1 ;
            rom[141] = 8'h43 ;
            rom[142] = 8'he3 ;
            rom[143] = 8'hde ;
            rom[144] = 8'hcd ;
            rom[145] = 8'hdc ;
            rom[146] = 8'h2f ;
            rom[147] = 8'hee ;
            rom[148] = 8'h30 ;
            rom[149] = 8'hed ;
            rom[150] = 8'hf6 ;
            rom[151] = 8'h97 ;
            rom[152] = 8'h18 ;
            rom[153] = 8'h25 ;
            rom[154] = 8'hd5 ;
            rom[155] = 8'h1c ;
            rom[156] = 8'h1e ;
            rom[157] = 8'hd9 ;
            rom[158] = 8'ha1 ;
            rom[159] = 8'h9f ;
            rom[160] = 8'h1f ;
            rom[161] = 8'hcd ;
            rom[162] = 8'h0e ;
            rom[163] = 8'h17 ;
            rom[164] = 8'hd1 ;
            rom[165] = 8'h19 ;
            rom[166] = 8'hed ;
            rom[167] = 8'hd4 ;
            rom[168] = 8'hc5 ;
            rom[169] = 8'h90 ;
            rom[170] = 8'h37 ;
            rom[171] = 8'h44 ;
            rom[172] = 8'he4 ;
            rom[173] = 8'hde ;
            rom[174] = 8'hdb ;
            rom[175] = 8'h29 ;
            rom[176] = 8'hc9 ;
            rom[177] = 8'hf6 ;
            rom[178] = 8'h39 ;
            rom[179] = 8'hbd ;
            rom[180] = 8'he4 ;
            rom[181] = 8'h4a ;
            rom[182] = 8'hfd ;
            rom[183] = 8'h21 ;
            rom[184] = 8'hf1 ;
            rom[185] = 8'h29 ;
            rom[186] = 8'hd8 ;
            rom[187] = 8'h3b ;
            rom[188] = 8'h58 ;
            rom[189] = 8'he3 ;
            rom[190] = 8'h19 ;
            rom[191] = 8'hb8 ;
            rom[192] = 8'h1e ;
            rom[193] = 8'h18 ;
            rom[194] = 8'hb9 ;
            rom[195] = 8'h24 ;
            rom[196] = 8'he0 ;
            rom[197] = 8'h21 ;
            rom[198] = 8'hcc ;
            rom[199] = 8'h9a ;
            rom[200] = 8'hdc ;
            rom[201] = 8'hbb ;
            rom[202] = 8'h29 ;
            rom[203] = 8'hf2 ;
            rom[204] = 8'h1d ;
            rom[205] = 8'h1b ;
            rom[206] = 8'hb6 ;
            rom[207] = 8'hfd ;
            rom[208] = 8'h43 ;
            rom[209] = 8'hd5 ;
            rom[210] = 8'hee ;
            rom[211] = 8'h00 ;
            rom[212] = 8'hca ;
            rom[213] = 8'ha0 ;
            rom[214] = 8'hdd ;
            rom[215] = 8'ha9 ;
            rom[216] = 8'hc6 ;
            rom[217] = 8'h04 ;
            rom[218] = 8'h81 ;
            rom[219] = 8'h04 ;
            rom[220] = 8'h2f ;
            rom[221] = 8'hed ;
            rom[222] = 8'h35 ;
            rom[223] = 8'h2e ;
            rom[224] = 8'h21 ;
            rom[225] = 8'h14 ;
            rom[226] = 8'hd3 ;
            rom[227] = 8'hb0 ;
            rom[228] = 8'h39 ;
            rom[229] = 8'hd5 ;
            rom[230] = 8'he1 ;
            rom[231] = 8'hc7 ;
            rom[232] = 8'hba ;
            rom[233] = 8'h15 ;
            rom[234] = 8'h1d ;
            rom[235] = 8'h1a ;
            rom[236] = 8'h1d ;
            rom[237] = 8'hc2 ;
            rom[238] = 8'hb2 ;
            rom[239] = 8'hb9 ;
            rom[240] = 8'h2c ;
            rom[241] = 8'h52 ;
            rom[242] = 8'h29 ;
            rom[243] = 8'hea ;
            rom[244] = 8'h4c ;
            rom[245] = 8'hf3 ;
            rom[246] = 8'hf4 ;
            rom[247] = 8'h47 ;
            rom[248] = 8'he5 ;
            rom[249] = 8'h3c ;
            rom[250] = 8'hf5 ;
            rom[251] = 8'hf8 ;
            rom[252] = 8'hfe ;
            rom[253] = 8'h33 ;
            rom[254] = 8'h42 ;
            rom[255] = 8'hf1 ;
            rom[256] = 8'h3e ;
            rom[257] = 8'h01 ;
            rom[258] = 8'hff ;
            rom[259] = 8'h57 ;
            rom[260] = 8'h2c ;
            rom[261] = 8'hee ;
            rom[262] = 8'h35 ;
            rom[263] = 8'hf0 ;
            rom[264] = 8'h38 ;
            rom[265] = 8'he6 ;
            rom[266] = 8'h38 ;
            rom[267] = 8'hd6 ;
            rom[268] = 8'h35 ;
            rom[269] = 8'he4 ;
            rom[270] = 8'hd7 ;
            rom[271] = 8'hb5 ;
            rom[272] = 8'h2d ;
            rom[273] = 8'hcd ;
            rom[274] = 8'h2e ;
            rom[275] = 8'h1c ;
            rom[276] = 8'hda ;
            rom[277] = 8'h28 ;
            rom[278] = 8'hcb ;
            rom[279] = 8'hc6 ;
            rom[280] = 8'h41 ;
            rom[281] = 8'h0c ;
            rom[282] = 8'hd3 ;
            rom[283] = 8'hdd ;
            rom[284] = 8'h4d ;
            rom[285] = 8'hdf ;
            rom[286] = 8'hd3 ;
            rom[287] = 8'hec ;
            rom[288] = 8'h3e ;
            rom[289] = 8'h27 ;
            rom[290] = 8'h16 ;
            rom[291] = 8'hc5 ;
            rom[292] = 8'hb6 ;
            rom[293] = 8'hd3 ;
            rom[294] = 8'h1b ;
            rom[295] = 8'h03 ;
            rom[296] = 8'hc5 ;
            rom[297] = 8'h17 ;
            rom[298] = 8'hb0 ;
            rom[299] = 8'h08 ;
            rom[300] = 8'h4c ;
            rom[301] = 8'h46 ;
            rom[302] = 8'hef ;
            rom[303] = 8'hc6 ;
            rom[304] = 8'hc8 ;
            rom[305] = 8'hd2 ;
            rom[306] = 8'hbd ;
            rom[307] = 8'hc3 ;
            rom[308] = 8'h01 ;
            rom[309] = 8'h42 ;
            rom[310] = 8'hf6 ;
            rom[311] = 8'hd6 ;
            rom[312] = 8'h2a ;
            rom[313] = 8'h3e ;
            rom[314] = 8'hd8 ;
            rom[315] = 8'h35 ;
            rom[316] = 8'h05 ;
            rom[317] = 8'h2d ;
            rom[318] = 8'heb ;
            rom[319] = 8'hb3 ;
            rom[320] = 8'hef ;
            rom[321] = 8'h02 ;
            rom[322] = 8'he9 ;
            rom[323] = 8'hcf ;
            rom[324] = 8'hd8 ;
            rom[325] = 8'hd4 ;
            rom[326] = 8'heb ;
            rom[327] = 8'he3 ;
            rom[328] = 8'h5e ;
            rom[329] = 8'h43 ;
            rom[330] = 8'h32 ;
            rom[331] = 8'hcd ;
            rom[332] = 8'h38 ;
            rom[333] = 8'h04 ;
            rom[334] = 8'h3c ;
            rom[335] = 8'hde ;
            rom[336] = 8'h3c ;
            rom[337] = 8'hcc ;
            rom[338] = 8'he7 ;
            rom[339] = 8'hf4 ;
            rom[340] = 8'hdf ;
            rom[341] = 8'hc1 ;
            rom[342] = 8'h3f ;
            rom[343] = 8'h2a ;
            rom[344] = 8'h4e ;
            rom[345] = 8'hff ;
            rom[346] = 8'h41 ;
            rom[347] = 8'hcb ;
            rom[348] = 8'had ;
            rom[349] = 8'hf5 ;
            rom[350] = 8'hcb ;
            rom[351] = 8'hd5 ;
            rom[352] = 8'hc6 ;
            rom[353] = 8'h32 ;
            rom[354] = 8'h35 ;
            rom[355] = 8'h3b ;
            rom[356] = 8'hcf ;
            rom[357] = 8'h2a ;
            rom[358] = 8'hd2 ;
            rom[359] = 8'h24 ;
            rom[360] = 8'hc7 ;
            rom[361] = 8'hba ;
            rom[362] = 8'h1e ;
            rom[363] = 8'h1f ;
            rom[364] = 8'hca ;
            rom[365] = 8'h17 ;
            rom[366] = 8'h29 ;
            rom[367] = 8'h04 ;
            rom[368] = 8'h2c ;
            rom[369] = 8'had ;
            rom[370] = 8'hde ;
            rom[371] = 8'hc5 ;
            rom[372] = 8'hd5 ;
            rom[373] = 8'h3b ;
            rom[374] = 8'h34 ;
            rom[375] = 8'h35 ;
            rom[376] = 8'hec ;
            rom[377] = 8'h3d ;
            rom[378] = 8'hcf ;
            rom[379] = 8'hc0 ;
            rom[380] = 8'h0b ;
            rom[381] = 8'ha0 ;
            rom[382] = 8'h24 ;
            rom[383] = 8'h13 ;
            rom[384] = 8'h1a ;
            rom[385] = 8'hbc ;
            rom[386] = 8'h18 ;
            rom[387] = 8'hbe ;
            rom[388] = 8'h42 ;
            rom[389] = 8'hb8 ;
            rom[390] = 8'hf8 ;
            rom[391] = 8'hef ;
            rom[392] = 8'hff ;
            rom[393] = 8'h04 ;
            rom[394] = 8'hfe ;
            rom[395] = 8'h49 ;
            rom[396] = 8'hed ;
            rom[397] = 8'h48 ;
            rom[398] = 8'hfc ;
            rom[399] = 8'h42 ;
            rom[400] = 8'hfb ;
            rom[401] = 8'h54 ;
            rom[402] = 8'hfa ;
            rom[403] = 8'heb ;
            rom[404] = 8'hf1 ;
            rom[405] = 8'hf5 ;
            rom[406] = 8'h69 ;
            rom[407] = 8'heb ;
            rom[408] = 8'h23 ;
            rom[409] = 8'h62 ;
            rom[410] = 8'hed ;
            rom[411] = 8'hf5 ;
            rom[412] = 8'hf6 ;
            rom[413] = 8'h27 ;
            rom[414] = 8'he4 ;
            rom[415] = 8'h43 ;
            rom[416] = 8'he3 ;
            rom[417] = 8'h53 ;
            rom[418] = 8'hf1 ;
            rom[419] = 8'h41 ;
            rom[420] = 8'h23 ;
            rom[421] = 8'hd6 ;
            rom[422] = 8'h2a ;
            rom[423] = 8'hde ;
            rom[424] = 8'h29 ;
            rom[425] = 8'hed ;
            rom[426] = 8'h1d ;
            rom[427] = 8'hcc ;
            rom[428] = 8'hc4 ;
            rom[429] = 8'h0e ;
            rom[430] = 8'h21 ;
            rom[431] = 8'h03 ;
            rom[432] = 8'h26 ;
            rom[433] = 8'hfd ;
            rom[434] = 8'hb4 ;
            rom[435] = 8'hce ;
            rom[436] = 8'h1d ;
            rom[437] = 8'hcd ;
            rom[438] = 8'hb1 ;
            rom[439] = 8'h25 ;
            rom[440] = 8'h0c ;
            rom[441] = 8'hca ;
            rom[442] = 8'hfa ;
            rom[443] = 8'h2f ;
            rom[444] = 8'h06 ;
            rom[445] = 8'hcf ;
            rom[446] = 8'h2e ;
            rom[447] = 8'hfc ;
            rom[448] = 8'h2b ;
            rom[449] = 8'hcc ;
            rom[450] = 8'h06 ;
            rom[451] = 8'hcd ;
            rom[452] = 8'h2e ;
            rom[453] = 8'hd7 ;
            rom[454] = 8'he9 ;
            rom[455] = 8'h36 ;
            rom[456] = 8'hd4 ;
            rom[457] = 8'h1d ;
            rom[458] = 8'hdf ;
            rom[459] = 8'hd0 ;
            rom[460] = 8'he5 ;
            rom[461] = 8'hd6 ;
            rom[462] = 8'hf8 ;
            rom[463] = 8'h31 ;
            rom[464] = 8'h2c ;
            rom[465] = 8'h37 ;
            rom[466] = 8'h44 ;
            rom[467] = 8'hca ;
            rom[468] = 8'hd0 ;
            rom[469] = 8'hcf ;
            rom[470] = 8'hbd ;
            rom[471] = 8'h02 ;
            rom[472] = 8'hd5 ;
            rom[473] = 8'h2c ;
            rom[474] = 8'hdf ;
            rom[475] = 8'hc3 ;
            rom[476] = 8'he3 ;
            rom[477] = 8'h09 ;
            rom[478] = 8'h2f ;
            rom[479] = 8'h29 ;
            rom[480] = 8'hb9 ;
            rom[481] = 8'hc7 ;
            rom[482] = 8'h35 ;
            rom[483] = 8'hf9 ;
            rom[484] = 8'h36 ;
            rom[485] = 8'h19 ;
            rom[486] = 8'h39 ;
            rom[487] = 8'h38 ;
            rom[488] = 8'hb3 ;
            rom[489] = 8'hc2 ;
            rom[490] = 8'he2 ;
            rom[491] = 8'h58 ;
            rom[492] = 8'he8 ;
            rom[493] = 8'hef ;
            rom[494] = 8'he4 ;
            rom[495] = 8'he4 ;
            rom[496] = 8'hd4 ;
            rom[497] = 8'he9 ;
            rom[498] = 8'h66 ;
            rom[499] = 8'h5a ;
            rom[500] = 8'h56 ;
            rom[501] = 8'h44 ;
            rom[502] = 8'he6 ;
            rom[503] = 8'hf1 ;
            rom[504] = 8'hd6 ;
            rom[505] = 8'h0a ;
            rom[506] = 8'h3a ;
            rom[507] = 8'hdb ;
            rom[508] = 8'h3f ;
            rom[509] = 8'hf6 ;
            rom[510] = 8'hcc ;
            rom[511] = 8'h42 ;
            rom[512] = 8'hdb ;
            rom[513] = 8'heb ;
            rom[514] = 8'h2d ;
            rom[515] = 8'hde ;
            rom[516] = 8'h33 ;
            rom[517] = 8'hda ;
            rom[518] = 8'h3e ;
            rom[519] = 8'h07 ;
            rom[520] = 8'h21 ;
            rom[521] = 8'h19 ;
            rom[522] = 8'h0a ;
            rom[523] = 8'hc3 ;
            rom[524] = 8'h1b ;
            rom[525] = 8'hc5 ;
            rom[526] = 8'hfe ;
            rom[527] = 8'ha2 ;
            rom[528] = 8'he7 ;
            rom[529] = 8'hc0 ;
            rom[530] = 8'h35 ;
            rom[531] = 8'hf0 ;
            rom[532] = 8'hea ;
            rom[533] = 8'hd7 ;
            rom[534] = 8'h1e ;
            rom[535] = 8'he5 ;
            rom[536] = 8'hfd ;
            rom[537] = 8'h43 ;
            rom[538] = 8'h51 ;
            rom[539] = 8'h0a ;
            rom[540] = 8'hf0 ;
            rom[541] = 8'hde ;
            rom[542] = 8'h21 ;
            rom[543] = 8'h1d ;
            rom[544] = 8'hd9 ;
            rom[545] = 8'hc8 ;
            rom[546] = 8'hf0 ;
            rom[547] = 8'h2c ;
            rom[548] = 8'h01 ;
            rom[549] = 8'h0f ;
            rom[550] = 8'ha6 ;
            rom[551] = 8'hc4 ;
            rom[552] = 8'h31 ;
            rom[553] = 8'h2f ;
            rom[554] = 8'h2d ;
            rom[555] = 8'h2d ;
            rom[556] = 8'h38 ;
            rom[557] = 8'hcd ;
            rom[558] = 8'hbe ;
            rom[559] = 8'heb ;
            rom[560] = 8'hf6 ;
            rom[561] = 8'hb0 ;
            rom[562] = 8'h04 ;
            rom[563] = 8'h38 ;
            rom[564] = 8'h4b ;
            rom[565] = 8'h44 ;
            rom[566] = 8'hd0 ;
            rom[567] = 8'h2f ;
            rom[568] = 8'h21 ;
            rom[569] = 8'h43 ;
            rom[570] = 8'he5 ;
            rom[571] = 8'hcc ;
            rom[572] = 8'hc7 ;
            rom[573] = 8'h26 ;
            rom[574] = 8'hdf ;
            rom[575] = 8'h2e ;
            rom[576] = 8'hc0 ;
            rom[577] = 8'h29 ;
            rom[578] = 8'h03 ;
            rom[579] = 8'h3e ;
            rom[580] = 8'h1c ;
            rom[581] = 8'h34 ;
            rom[582] = 8'h2d ;
            rom[583] = 8'hdc ;
            rom[584] = 8'hb1 ;
            rom[585] = 8'hd8 ;
            rom[586] = 8'hc8 ;
            rom[587] = 8'h2a ;
            rom[588] = 8'hfd ;
            rom[589] = 8'h37 ;
            rom[590] = 8'h32 ;
            rom[591] = 8'h45 ;
            rom[592] = 8'hff ;
            rom[593] = 8'h30 ;
            rom[594] = 8'h1b ;
            rom[595] = 8'h35 ;
            rom[596] = 8'hc3 ;
            rom[597] = 8'hb0 ;
            rom[598] = 8'hc7 ;
            rom[599] = 8'h44 ;
            rom[600] = 8'h27 ;
            rom[601] = 8'h2a ;
            rom[602] = 8'hfe ;
            rom[603] = 8'hf8 ;
            rom[604] = 8'hd8 ;
            rom[605] = 8'h06 ;
            rom[606] = 8'h31 ;
            rom[607] = 8'h4d ;
            rom[608] = 8'h3a ;
            rom[609] = 8'he9 ;
            rom[610] = 8'h21 ;
            rom[611] = 8'h28 ;
            rom[612] = 8'hc5 ;
            rom[613] = 8'he2 ;
            rom[614] = 8'hb6 ;
            rom[615] = 8'h1c ;
            rom[616] = 8'hd2 ;
            rom[617] = 8'h1b ;
            rom[618] = 8'hb8 ;
            rom[619] = 8'h22 ;
            rom[620] = 8'hdf ;
            rom[621] = 8'hd2 ;
            rom[622] = 8'h31 ;
            rom[623] = 8'hf9 ;
            rom[624] = 8'h1a ;
            rom[625] = 8'h3b ;
            rom[626] = 8'h32 ;
            rom[627] = 8'hdc ;
            rom[628] = 8'h3e ;
            rom[629] = 8'hde ;
            rom[630] = 8'h15 ;
            rom[631] = 8'h01 ;
            rom[632] = 8'hd0 ;
            rom[633] = 8'hc2 ;
            rom[634] = 8'hba ;
            rom[635] = 8'hba ;
            rom[636] = 8'hbb ;
            rom[637] = 8'h19 ;
            rom[638] = 8'hb8 ;
            rom[639] = 8'h07 ;
            rom[640] = 8'h2f ;
            rom[641] = 8'hc2 ;
            rom[642] = 8'h23 ;
            rom[643] = 8'h1b ;
            rom[644] = 8'h32 ;
            rom[645] = 8'h0d ;
            rom[646] = 8'hca ;
            rom[647] = 8'hc5 ;
            rom[648] = 8'hfa ;
            rom[649] = 8'hed ;
            rom[650] = 8'he5 ;
            rom[651] = 8'h17 ;
            rom[652] = 8'h28 ;
            rom[653] = 8'hec ;
            rom[654] = 8'h2c ;
            rom[655] = 8'hc3 ;
            rom[656] = 8'h0c ;
            rom[657] = 8'hd6 ;
            rom[658] = 8'he1 ;
            rom[659] = 8'h00 ;
            rom[660] = 8'hf8 ;
            rom[661] = 8'h44 ;
            rom[662] = 8'h53 ;
            rom[663] = 8'he1 ;
            rom[664] = 8'hd7 ;
            rom[665] = 8'h02 ;
            rom[666] = 8'h40 ;
            rom[667] = 8'he0 ;
            rom[668] = 8'hfa ;
            rom[669] = 8'h4a ;
            rom[670] = 8'he2 ;
            rom[671] = 8'h61 ;
            rom[672] = 8'hf9 ;
            rom[673] = 8'hee ;
            rom[674] = 8'he4 ;
            rom[675] = 8'he4 ;
            rom[676] = 8'hfb ;
            rom[677] = 8'hd7 ;
            rom[678] = 8'he3 ;
            rom[679] = 8'h61 ;
            rom[680] = 8'h0c ;
            rom[681] = 8'hc1 ;
            rom[682] = 8'h0b ;
            rom[683] = 8'h1c ;
            rom[684] = 8'hcf ;
            rom[685] = 8'h20 ;
            rom[686] = 8'h16 ;
            rom[687] = 8'hd2 ;
            rom[688] = 8'hc0 ;
            rom[689] = 8'hd5 ;
            rom[690] = 8'he3 ;
            rom[691] = 8'h47 ;
            rom[692] = 8'hdf ;
            rom[693] = 8'hec ;
            rom[694] = 8'hdc ;
            rom[695] = 8'hd6 ;
            rom[696] = 8'hd8 ;
            rom[697] = 8'hde ;
            rom[698] = 8'hd2 ;
            rom[699] = 8'h3f ;
            rom[700] = 8'hec ;
            rom[701] = 8'h3c ;
            rom[702] = 8'hc9 ;
            rom[703] = 8'h03 ;
            rom[704] = 8'h35 ;
            rom[705] = 8'he8 ;
            rom[706] = 8'hba ;
            rom[707] = 8'hd9 ;
            rom[708] = 8'h26 ;
            rom[709] = 8'hea ;
            rom[710] = 8'h01 ;
            rom[711] = 8'h47 ;
            rom[712] = 8'h3d ;
            rom[713] = 8'h11 ;
            rom[714] = 8'he3 ;
            rom[715] = 8'h40 ;
            rom[716] = 8'h36 ;
            rom[717] = 8'hf0 ;
            rom[718] = 8'hf8 ;
            rom[719] = 8'hf2 ;
            rom[720] = 8'hdc ;
            rom[721] = 8'hfc ;
            rom[722] = 8'h25 ;
            rom[723] = 8'h0c ;
            rom[724] = 8'h32 ;
            rom[725] = 8'h40 ;
            rom[726] = 8'hd9 ;
            rom[727] = 8'h49 ;
            rom[728] = 8'hd5 ;
            rom[729] = 8'h1f ;
            rom[730] = 8'hbb ;
            rom[731] = 8'hce ;
            rom[732] = 8'h26 ;
            rom[733] = 8'h25 ;
            rom[734] = 8'hd4 ;
            rom[735] = 8'h13 ;
            rom[736] = 8'h34 ;
            rom[737] = 8'h2b ;
            rom[738] = 8'hcd ;
            rom[739] = 8'hbd ;
            rom[740] = 8'h02 ;
            rom[741] = 8'h2c ;
            rom[742] = 8'hdd ;
            rom[743] = 8'he0 ;
            rom[744] = 8'h4e ;
            rom[745] = 8'hd7 ;
            rom[746] = 8'hef ;
            rom[747] = 8'h29 ;
            rom[748] = 8'hd6 ;
            rom[749] = 8'h15 ;
            rom[750] = 8'hb9 ;
            rom[751] = 8'hbb ;
            rom[752] = 8'h0e ;
            rom[753] = 8'hfe ;
            rom[754] = 8'hd0 ;
            rom[755] = 8'hc8 ;
            rom[756] = 8'h13 ;
            rom[757] = 8'h1f ;
            rom[758] = 8'h17 ;
            rom[759] = 8'hde ;
            rom[760] = 8'hfe ;
            rom[761] = 8'h02 ;
            rom[762] = 8'h2d ;
            rom[763] = 8'hda ;
            rom[764] = 8'hd8 ;
            rom[765] = 8'h08 ;
            rom[766] = 8'h13 ;
            rom[767] = 8'hd9 ;
            rom[768] = 8'h10 ;
            rom[769] = 8'hf1 ;
            rom[770] = 8'h3e ;
            rom[771] = 8'h47 ;
            rom[772] = 8'hea ;
            rom[773] = 8'hdb ;
            rom[774] = 8'hd0 ;
            rom[775] = 8'he0 ;
            rom[776] = 8'hc5 ;
            rom[777] = 8'h58 ;
            rom[778] = 8'h4d ;
            rom[779] = 8'h4d ;
            rom[780] = 8'h08 ;
            rom[781] = 8'h44 ;
            rom[782] = 8'h40 ;
            rom[783] = 8'he5 ;
            rom[784] = 8'h27 ;
            rom[785] = 8'hda ;
            rom[786] = 8'h3c ;
            rom[787] = 8'h2f ;
            rom[788] = 8'hdb ;
            rom[789] = 8'hed ;
            rom[790] = 8'hcd ;
            rom[791] = 8'hfa ;
            rom[792] = 8'hc8 ;
            rom[793] = 8'h1e ;
            rom[794] = 8'hdd ;
            rom[795] = 8'hda ;
            rom[796] = 8'h24 ;
            rom[797] = 8'he9 ;
            rom[798] = 8'h13 ;
            rom[799] = 8'he2 ;
            rom[800] = 8'h21 ;
            rom[801] = 8'he8 ;
            rom[802] = 8'h25 ;
            rom[803] = 8'h05 ;
            rom[804] = 8'hcc ;
            rom[805] = 8'hde ;
            rom[806] = 8'h33 ;
            rom[807] = 8'hc4 ;
            rom[808] = 8'hc2 ;
            rom[809] = 8'hfd ;
            rom[810] = 8'hcd ;
            rom[811] = 8'h3e ;
            rom[812] = 8'h34 ;
            rom[813] = 8'h19 ;
            rom[814] = 8'hf1 ;
            rom[815] = 8'hfe ;
            rom[816] = 8'he6 ;
            rom[817] = 8'hb7 ;
            rom[818] = 8'hec ;
            rom[819] = 8'h41 ;
            rom[820] = 8'hdb ;
            rom[821] = 8'hda ;
            rom[822] = 8'hcf ;
            rom[823] = 8'h06 ;
            rom[824] = 8'h1f ;
            rom[825] = 8'h24 ;
            rom[826] = 8'h3a ;
            rom[827] = 8'h2f ;
            rom[828] = 8'hca ;
            rom[829] = 8'hc1 ;
            rom[830] = 8'he4 ;
            rom[831] = 8'hcd ;
            rom[832] = 8'h3b ;
            rom[833] = 8'he9 ;
            rom[834] = 8'h2c ;
            rom[835] = 8'h37 ;
            rom[836] = 8'h3c ;
            rom[837] = 8'he2 ;
            rom[838] = 8'he0 ;
            rom[839] = 8'he9 ;
            rom[840] = 8'hcd ;
            rom[841] = 8'h39 ;
            rom[842] = 8'he1 ;
            rom[843] = 8'hdb ;
            rom[844] = 8'hce ;
            rom[845] = 8'hd2 ;
            rom[846] = 8'h2e ;
            rom[847] = 8'hc4 ;
            rom[848] = 8'hdc ;
            rom[849] = 8'h49 ;
            rom[850] = 8'hda ;
            rom[851] = 8'h1d ;
            rom[852] = 8'hc7 ;
            rom[853] = 8'h2a ;
            rom[854] = 8'hce ;
            rom[855] = 8'hee ;
            rom[856] = 8'hca ;
            rom[857] = 8'hc0 ;
            rom[858] = 8'heb ;
            rom[859] = 8'hd3 ;
            rom[860] = 8'hea ;
            rom[861] = 8'h3d ;
            rom[862] = 8'hec ;
            rom[863] = 8'hdb ;
            rom[864] = 8'h39 ;
            rom[865] = 8'he7 ;
            rom[866] = 8'h22 ;
            rom[867] = 8'he1 ;
            rom[868] = 8'h10 ;
            rom[869] = 8'hfc ;
            rom[870] = 8'hbf ;
            rom[871] = 8'h87 ;
            rom[872] = 8'h92 ;
            rom[873] = 8'hf1 ;
            rom[874] = 8'hef ;
            rom[875] = 8'h3f ;
            rom[876] = 8'h15 ;
            rom[877] = 8'hfe ;
            rom[878] = 8'hd2 ;
            rom[879] = 8'hbe ;
            rom[880] = 8'hd9 ;
            rom[881] = 8'hf0 ;
            rom[882] = 8'he8 ;
            rom[883] = 8'hcd ;
            rom[884] = 8'hd9 ;
            rom[885] = 8'heb ;
            rom[886] = 8'hdc ;
            rom[887] = 8'he7 ;
            rom[888] = 8'h4e ;
            rom[889] = 8'h3f ;
            rom[890] = 8'h51 ;
            rom[891] = 8'h7b ;
            rom[892] = 8'h15 ;
            rom[893] = 8'h2d ;
            rom[894] = 8'h65 ;
            rom[895] = 8'h77 ;
            rom[896] = 8'hf8 ;
            rom[897] = 8'hdd ;
            rom[898] = 8'h49 ;
            rom[899] = 8'h58 ;
            rom[900] = 8'he1 ;
            rom[901] = 8'hcd ;
            rom[902] = 8'hcb ;
            rom[903] = 8'hec ;
            rom[904] = 8'hf0 ;
            rom[905] = 8'hd7 ;
            rom[906] = 8'h26 ;
            rom[907] = 8'h29 ;
            rom[908] = 8'hc5 ;
            rom[909] = 8'h12 ;
            rom[910] = 8'hd8 ;
            rom[911] = 8'h45 ;
            rom[912] = 8'h4e ;
            rom[913] = 8'h27 ;
            rom[914] = 8'h1b ;
            rom[915] = 8'h69 ;
            rom[916] = 8'h75 ;
            rom[917] = 8'h5a ;
            rom[918] = 8'h63 ;
            rom[919] = 8'h32 ;
            rom[920] = 8'h1c ;
            rom[921] = 8'ha3 ;
            rom[922] = 8'h25 ;
            rom[923] = 8'h22 ;
            rom[924] = 8'h2a ;
            rom[925] = 8'h73 ;
            rom[926] = 8'h91 ;
            rom[927] = 8'h17 ;
            rom[928] = 8'h70 ;
            rom[929] = 8'h79 ;
            rom[930] = 8'h27 ;
            rom[931] = 8'h32 ;
            rom[932] = 8'h16 ;
            rom[933] = 8'hd5 ;
            rom[934] = 8'h66 ;
            rom[935] = 8'hbf ;
            rom[936] = 8'hd3 ;
            rom[937] = 8'haa ;
            rom[938] = 8'h2c ;
            rom[939] = 8'hce ;
            rom[940] = 8'h31 ;
            rom[941] = 8'he3 ;
            rom[942] = 8'hdc ;
            rom[943] = 8'he8 ;
            rom[944] = 8'h39 ;
            rom[945] = 8'hed ;
            rom[946] = 8'hfe ;
            rom[947] = 8'h43 ;
            rom[948] = 8'h24 ;
            rom[949] = 8'hc1 ;
            rom[950] = 8'h39 ;
            rom[951] = 8'h05 ;
            rom[952] = 8'hf8 ;
            rom[953] = 8'hee ;
            rom[954] = 8'h35 ;
            rom[955] = 8'h04 ;
            rom[956] = 8'hda ;
            rom[957] = 8'h27 ;
            rom[958] = 8'hce ;
            rom[959] = 8'hc2 ;
            rom[960] = 8'h0d ;
            rom[961] = 8'hac ;
            rom[962] = 8'hb5 ;
            rom[963] = 8'h22 ;
            rom[964] = 8'hc6 ;
            rom[965] = 8'hf3 ;
            rom[966] = 8'hac ;
            rom[967] = 8'h0e ;
            rom[968] = 8'h14 ;
            rom[969] = 8'hd2 ;
            rom[970] = 8'h34 ;
            rom[971] = 8'hde ;
            rom[972] = 8'h35 ;
            rom[973] = 8'hda ;
            rom[974] = 8'hca ;
            rom[975] = 8'hdf ;
            rom[976] = 8'h2e ;
            rom[977] = 8'hd5 ;
            rom[978] = 8'h3b ;
            rom[979] = 8'he5 ;
            rom[980] = 8'h4b ;
            rom[981] = 8'h52 ;
            rom[982] = 8'hd8 ;
            rom[983] = 8'he1 ;
            rom[984] = 8'hd2 ;
            rom[985] = 8'hd8 ;
            rom[986] = 8'hd4 ;
            rom[987] = 8'hc4 ;
            rom[988] = 8'h4e ;
            rom[989] = 8'h5a ;
            rom[990] = 8'hb0 ;
            rom[991] = 8'h00 ;
            rom[992] = 8'h10 ;
            rom[993] = 8'hc0 ;
            rom[994] = 8'h15 ;
            rom[995] = 8'h07 ;
            rom[996] = 8'hf4 ;
            rom[997] = 8'h19 ;
            rom[998] = 8'haf ;
            rom[999] = 8'haa ;
            rom[1000] = 8'hc9 ;
            rom[1001] = 8'h52 ;
            rom[1002] = 8'hf0 ;
            rom[1003] = 8'hd6 ;
            rom[1004] = 8'he7 ;
            rom[1005] = 8'hdc ;
            rom[1006] = 8'hf3 ;
            rom[1007] = 8'h08 ;
            rom[1008] = 8'h5c ;
            rom[1009] = 8'h58 ;
            rom[1010] = 8'h4e ;
            rom[1011] = 8'h4e ;
            rom[1012] = 8'hd4 ;
            rom[1013] = 8'hd5 ;
            rom[1014] = 8'hd9 ;
            rom[1015] = 8'hc5 ;
            rom[1016] = 8'he7 ;
            rom[1017] = 8'hc7 ;
            rom[1018] = 8'h59 ;
            rom[1019] = 8'h52 ;
            rom[1020] = 8'hae ;
            rom[1021] = 8'hca ;
            rom[1022] = 8'h14 ;
            rom[1023] = 8'hdd ;
            rom[1024] = 8'hbd ;
            rom[1025] = 8'h0c ;
            rom[1026] = 8'h0e ;
            rom[1027] = 8'h1f ;
            rom[1028] = 8'hca ;
            rom[1029] = 8'h2c ;
            rom[1030] = 8'he4 ;
            rom[1031] = 8'he7 ;
            rom[1032] = 8'hed ;
            rom[1033] = 8'hff ;
            rom[1034] = 8'h3d ;
            rom[1035] = 8'hfd ;
            rom[1036] = 8'h0a ;
            rom[1037] = 8'h46 ;
            rom[1038] = 8'h14 ;
            rom[1039] = 8'he9 ;
            rom[1040] = 8'hdf ;
            rom[1041] = 8'h2d ;
            rom[1042] = 8'hd7 ;
            rom[1043] = 8'hd3 ;
            rom[1044] = 8'hfb ;
            rom[1045] = 8'h16 ;
            rom[1046] = 8'he1 ;
            rom[1047] = 8'hce ;
            rom[1048] = 8'h57 ;
            rom[1049] = 8'hcb ;
            rom[1050] = 8'h2b ;
            rom[1051] = 8'hb7 ;
            rom[1052] = 8'h39 ;
            rom[1053] = 8'hf2 ;
            rom[1054] = 8'h29 ;
            rom[1055] = 8'hd1 ;
            rom[1056] = 8'hf3 ;
            rom[1057] = 8'he0 ;
            rom[1058] = 8'h34 ;
            rom[1059] = 8'he4 ;
            rom[1060] = 8'h0c ;
            rom[1061] = 8'hae ;
            rom[1062] = 8'he4 ;
            rom[1063] = 8'he9 ;
            rom[1064] = 8'h21 ;
            rom[1065] = 8'h11 ;
            rom[1066] = 8'hca ;
            rom[1067] = 8'hd3 ;
            rom[1068] = 8'h33 ;
            rom[1069] = 8'hb1 ;
            rom[1070] = 8'hdc ;
            rom[1071] = 8'hfd ;
            rom[1072] = 8'hdc ;
            rom[1073] = 8'hf0 ;
            rom[1074] = 8'h1c ;
            rom[1075] = 8'h29 ;
            rom[1076] = 8'h53 ;
            rom[1077] = 8'h33 ;
            rom[1078] = 8'hfa ;
            rom[1079] = 8'hd9 ;
            rom[1080] = 8'h02 ;
            rom[1081] = 8'h21 ;
            rom[1082] = 8'hf0 ;
            rom[1083] = 8'h1a ;
            rom[1084] = 8'hc6 ;
            rom[1085] = 8'hfb ;
            rom[1086] = 8'ha9 ;
            rom[1087] = 8'hc9 ;
            rom[1088] = 8'h04 ;
            rom[1089] = 8'hf7 ;
            rom[1090] = 8'he0 ;
            rom[1091] = 8'h50 ;
            rom[1092] = 8'h37 ;
            rom[1093] = 8'h46 ;
            rom[1094] = 8'hed ;
            rom[1095] = 8'h06 ;
            rom[1096] = 8'h42 ;
            rom[1097] = 8'h07 ;
            rom[1098] = 8'hec ;
            rom[1099] = 8'hc2 ;
            rom[1100] = 8'heb ;
            rom[1101] = 8'hc9 ;
            rom[1102] = 8'h13 ;
            rom[1103] = 8'hd3 ;
            rom[1104] = 8'hc5 ;
            rom[1105] = 8'h14 ;
            rom[1106] = 8'hce ;
            rom[1107] = 8'h0c ;
            rom[1108] = 8'h37 ;
            rom[1109] = 8'h34 ;
            rom[1110] = 8'hde ;
            rom[1111] = 8'h35 ;
            rom[1112] = 8'he8 ;
            rom[1113] = 8'h3d ;
            rom[1114] = 8'he0 ;
            rom[1115] = 8'h21 ;
            rom[1116] = 8'he3 ;
            rom[1117] = 8'h36 ;
            rom[1118] = 8'hc1 ;
            rom[1119] = 8'h2d ;
            rom[1120] = 8'h3d ;
            rom[1121] = 8'h2d ;
            rom[1122] = 8'hcd ;
            rom[1123] = 8'h01 ;
            rom[1124] = 8'hcb ;
            rom[1125] = 8'hdd ;
            rom[1126] = 8'h49 ;
            rom[1127] = 8'hd2 ;
            rom[1128] = 8'h0e ;
            rom[1129] = 8'h38 ;
            rom[1130] = 8'hc5 ;
            rom[1131] = 8'h44 ;
            rom[1132] = 8'hf2 ;
            rom[1133] = 8'hea ;
            rom[1134] = 8'hf2 ;
            rom[1135] = 8'h23 ;
            rom[1136] = 8'h22 ;
            rom[1137] = 8'hdc ;
            rom[1138] = 8'hd9 ;
            rom[1139] = 8'h44 ;
            rom[1140] = 8'h32 ;
            rom[1141] = 8'h1d ;
            rom[1142] = 8'hda ;
            rom[1143] = 8'hee ;
            rom[1144] = 8'h2b ;
            rom[1145] = 8'hc7 ;
            rom[1146] = 8'hdd ;
            rom[1147] = 8'hba ;
            rom[1148] = 8'hba ;
            rom[1149] = 8'h2f ;
            rom[1150] = 8'he4 ;
            rom[1151] = 8'hdb ;
        end
    always
        @(*)
        begin
            data <=  rom[addr] ;
        end
endmodule



