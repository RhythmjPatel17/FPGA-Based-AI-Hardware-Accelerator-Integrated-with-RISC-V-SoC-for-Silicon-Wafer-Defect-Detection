(* keep_hierarchy = "yes", dont_touch = "true" *)

module weights_rom_1 (
    input wire [9:0] addr, 
    output reg [7:0] data) ;
    reg [7:0] rom [0:863] ; 
    initial
        begin
            rom[0] = 8'h20 ;
            rom[1] = 8'h02 ;
            rom[2] = 8'hc2 ;
            rom[3] = 8'h33 ;
            rom[4] = 8'he7 ;
            rom[5] = 8'h29 ;
            rom[6] = 8'hca ;
            rom[7] = 8'h2b ;
            rom[8] = 8'hd8 ;
            rom[9] = 8'h83 ;
            rom[10] = 8'h41 ;
            rom[11] = 8'hdf ;
            rom[12] = 8'hee ;
            rom[13] = 8'hef ;
            rom[14] = 8'hdd ;
            rom[15] = 8'h41 ;
            rom[16] = 8'h03 ;
            rom[17] = 8'h3b ;
            rom[18] = 8'hbd ;
            rom[19] = 8'h17 ;
            rom[20] = 8'haf ;
            rom[21] = 8'h2f ;
            rom[22] = 8'he3 ;
            rom[23] = 8'hfa ;
            rom[24] = 8'hd7 ;
            rom[25] = 8'h22 ;
            rom[26] = 8'he9 ;
            rom[27] = 8'h3a ;
            rom[28] = 8'h2e ;
            rom[29] = 8'hf4 ;
            rom[30] = 8'he0 ;
            rom[31] = 8'hde ;
            rom[32] = 8'hfc ;
            rom[33] = 8'hf8 ;
            rom[34] = 8'h0f ;
            rom[35] = 8'h04 ;
            rom[36] = 8'he6 ;
            rom[37] = 8'hf6 ;
            rom[38] = 8'hdd ;
            rom[39] = 8'hf1 ;
            rom[40] = 8'h17 ;
            rom[41] = 8'ha8 ;
            rom[42] = 8'h42 ;
            rom[43] = 8'hdf ;
            rom[44] = 8'h09 ;
            rom[45] = 8'h26 ;
            rom[46] = 8'hfa ;
            rom[47] = 8'he4 ;
            rom[48] = 8'h02 ;
            rom[49] = 8'h18 ;
            rom[50] = 8'hf0 ;
            rom[51] = 8'hf4 ;
            rom[52] = 8'hb8 ;
            rom[53] = 8'h51 ;
            rom[54] = 8'hde ;
            rom[55] = 8'h43 ;
            rom[56] = 8'hf4 ;
            rom[57] = 8'hee ;
            rom[58] = 8'h2e ;
            rom[59] = 8'h07 ;
            rom[60] = 8'hc4 ;
            rom[61] = 8'h19 ;
            rom[62] = 8'hb7 ;
            rom[63] = 8'h2b ;
            rom[64] = 8'hbe ;
            rom[65] = 8'hf3 ;
            rom[66] = 8'hd6 ;
            rom[67] = 8'hf9 ;
            rom[68] = 8'hcb ;
            rom[69] = 8'h08 ;
            rom[70] = 8'hf7 ;
            rom[71] = 8'h16 ;
            rom[72] = 8'h14 ;
            rom[73] = 8'h81 ;
            rom[74] = 8'h34 ;
            rom[75] = 8'he4 ;
            rom[76] = 8'hc3 ;
            rom[77] = 8'hdc ;
            rom[78] = 8'he7 ;
            rom[79] = 8'hea ;
            rom[80] = 8'hc6 ;
            rom[81] = 8'h4c ;
            rom[82] = 8'hd7 ;
            rom[83] = 8'hf2 ;
            rom[84] = 8'heb ;
            rom[85] = 8'h17 ;
            rom[86] = 8'hcd ;
            rom[87] = 8'h11 ;
            rom[88] = 8'h23 ;
            rom[89] = 8'hf5 ;
            rom[90] = 8'h08 ;
            rom[91] = 8'h29 ;
            rom[92] = 8'hdc ;
            rom[93] = 8'h0d ;
            rom[94] = 8'hc8 ;
            rom[95] = 8'hf5 ;
            rom[96] = 8'h07 ;
            rom[97] = 8'h13 ;
            rom[98] = 8'he5 ;
            rom[99] = 8'h19 ;
            rom[100] = 8'h24 ;
            rom[101] = 8'h43 ;
            rom[102] = 8'hb8 ;
            rom[103] = 8'h53 ;
            rom[104] = 8'he6 ;
            rom[105] = 8'h1a ;
            rom[106] = 8'h20 ;
            rom[107] = 8'hdd ;
            rom[108] = 8'hea ;
            rom[109] = 8'hdf ;
            rom[110] = 8'hc2 ;
            rom[111] = 8'hee ;
            rom[112] = 8'h2d ;
            rom[113] = 8'hc6 ;
            rom[114] = 8'hd8 ;
            rom[115] = 8'h18 ;
            rom[116] = 8'h1f ;
            rom[117] = 8'hfb ;
            rom[118] = 8'he4 ;
            rom[119] = 8'ha7 ;
            rom[120] = 8'hbd ;
            rom[121] = 8'h22 ;
            rom[122] = 8'h20 ;
            rom[123] = 8'h2c ;
            rom[124] = 8'h1d ;
            rom[125] = 8'hac ;
            rom[126] = 8'hcf ;
            rom[127] = 8'h14 ;
            rom[128] = 8'hf4 ;
            rom[129] = 8'hed ;
            rom[130] = 8'he4 ;
            rom[131] = 8'h02 ;
            rom[132] = 8'hd3 ;
            rom[133] = 8'h5f ;
            rom[134] = 8'hc6 ;
            rom[135] = 8'hfd ;
            rom[136] = 8'hf9 ;
            rom[137] = 8'he0 ;
            rom[138] = 8'hef ;
            rom[139] = 8'h26 ;
            rom[140] = 8'hcc ;
            rom[141] = 8'h28 ;
            rom[142] = 8'hee ;
            rom[143] = 8'hdb ;
            rom[144] = 8'hff ;
            rom[145] = 8'h9d ;
            rom[146] = 8'h15 ;
            rom[147] = 8'h10 ;
            rom[148] = 8'hd6 ;
            rom[149] = 8'hd9 ;
            rom[150] = 8'hb1 ;
            rom[151] = 8'hef ;
            rom[152] = 8'hf0 ;
            rom[153] = 8'heb ;
            rom[154] = 8'h2a ;
            rom[155] = 8'hf6 ;
            rom[156] = 8'hc8 ;
            rom[157] = 8'he6 ;
            rom[158] = 8'hd8 ;
            rom[159] = 8'h2f ;
            rom[160] = 8'heb ;
            rom[161] = 8'hd8 ;
            rom[162] = 8'hff ;
            rom[163] = 8'hbd ;
            rom[164] = 8'hce ;
            rom[165] = 8'h50 ;
            rom[166] = 8'hdf ;
            rom[167] = 8'hd4 ;
            rom[168] = 8'hda ;
            rom[169] = 8'hf1 ;
            rom[170] = 8'h03 ;
            rom[171] = 8'he2 ;
            rom[172] = 8'hfc ;
            rom[173] = 8'h3c ;
            rom[174] = 8'hf8 ;
            rom[175] = 8'h0f ;
            rom[176] = 8'hc7 ;
            rom[177] = 8'hb7 ;
            rom[178] = 8'h14 ;
            rom[179] = 8'hec ;
            rom[180] = 8'hfe ;
            rom[181] = 8'h07 ;
            rom[182] = 8'ha0 ;
            rom[183] = 8'h9e ;
            rom[184] = 8'h1a ;
            rom[185] = 8'hf5 ;
            rom[186] = 8'hf8 ;
            rom[187] = 8'h19 ;
            rom[188] = 8'hfa ;
            rom[189] = 8'h1a ;
            rom[190] = 8'he6 ;
            rom[191] = 8'h29 ;
            rom[192] = 8'h2a ;
            rom[193] = 8'hd5 ;
            rom[194] = 8'h4f ;
            rom[195] = 8'h03 ;
            rom[196] = 8'h38 ;
            rom[197] = 8'he9 ;
            rom[198] = 8'hee ;
            rom[199] = 8'h07 ;
            rom[200] = 8'he5 ;
            rom[201] = 8'hf7 ;
            rom[202] = 8'hb7 ;
            rom[203] = 8'hea ;
            rom[204] = 8'he4 ;
            rom[205] = 8'hee ;
            rom[206] = 8'hcd ;
            rom[207] = 8'h08 ;
            rom[208] = 8'hd0 ;
            rom[209] = 8'h3a ;
            rom[210] = 8'hdd ;
            rom[211] = 8'h31 ;
            rom[212] = 8'h31 ;
            rom[213] = 8'hfb ;
            rom[214] = 8'hf3 ;
            rom[215] = 8'haa ;
            rom[216] = 8'hdb ;
            rom[217] = 8'h26 ;
            rom[218] = 8'h10 ;
            rom[219] = 8'h4d ;
            rom[220] = 8'h27 ;
            rom[221] = 8'hbc ;
            rom[222] = 8'hfe ;
            rom[223] = 8'h13 ;
            rom[224] = 8'h1d ;
            rom[225] = 8'h03 ;
            rom[226] = 8'hff ;
            rom[227] = 8'hea ;
            rom[228] = 8'h3d ;
            rom[229] = 8'he3 ;
            rom[230] = 8'hf2 ;
            rom[231] = 8'hc0 ;
            rom[232] = 8'h17 ;
            rom[233] = 8'he7 ;
            rom[234] = 8'hb0 ;
            rom[235] = 8'h0a ;
            rom[236] = 8'hf7 ;
            rom[237] = 8'he9 ;
            rom[238] = 8'hd5 ;
            rom[239] = 8'h0f ;
            rom[240] = 8'hdd ;
            rom[241] = 8'h14 ;
            rom[242] = 8'he7 ;
            rom[243] = 8'h2a ;
            rom[244] = 8'he2 ;
            rom[245] = 8'hff ;
            rom[246] = 8'h23 ;
            rom[247] = 8'h0f ;
            rom[248] = 8'hd4 ;
            rom[249] = 8'hdf ;
            rom[250] = 8'hcd ;
            rom[251] = 8'h16 ;
            rom[252] = 8'he6 ;
            rom[253] = 8'hfe ;
            rom[254] = 8'h3c ;
            rom[255] = 8'h30 ;
            rom[256] = 8'hfa ;
            rom[257] = 8'h0b ;
            rom[258] = 8'h07 ;
            rom[259] = 8'h22 ;
            rom[260] = 8'h06 ;
            rom[261] = 8'hf6 ;
            rom[262] = 8'h46 ;
            rom[263] = 8'ha0 ;
            rom[264] = 8'hea ;
            rom[265] = 8'hd5 ;
            rom[266] = 8'hd3 ;
            rom[267] = 8'h1d ;
            rom[268] = 8'hdb ;
            rom[269] = 8'h1a ;
            rom[270] = 8'hdb ;
            rom[271] = 8'hc7 ;
            rom[272] = 8'h16 ;
            rom[273] = 8'he5 ;
            rom[274] = 8'hd0 ;
            rom[275] = 8'he6 ;
            rom[276] = 8'hcb ;
            rom[277] = 8'hdc ;
            rom[278] = 8'hfe ;
            rom[279] = 8'hdc ;
            rom[280] = 8'h30 ;
            rom[281] = 8'h0e ;
            rom[282] = 8'hdb ;
            rom[283] = 8'h31 ;
            rom[284] = 8'h2b ;
            rom[285] = 8'h3d ;
            rom[286] = 8'h3b ;
            rom[287] = 8'hcb ;
            rom[288] = 8'h56 ;
            rom[289] = 8'he7 ;
            rom[290] = 8'h1a ;
            rom[291] = 8'hea ;
            rom[292] = 8'h02 ;
            rom[293] = 8'hf4 ;
            rom[294] = 8'hd2 ;
            rom[295] = 8'hc1 ;
            rom[296] = 8'he4 ;
            rom[297] = 8'hc9 ;
            rom[298] = 8'h33 ;
            rom[299] = 8'h1f ;
            rom[300] = 8'h17 ;
            rom[301] = 8'heb ;
            rom[302] = 8'hd1 ;
            rom[303] = 8'h3f ;
            rom[304] = 8'h54 ;
            rom[305] = 8'h12 ;
            rom[306] = 8'hfa ;
            rom[307] = 8'hde ;
            rom[308] = 8'haf ;
            rom[309] = 8'h0b ;
            rom[310] = 8'h3b ;
            rom[311] = 8'h2e ;
            rom[312] = 8'h31 ;
            rom[313] = 8'he1 ;
            rom[314] = 8'h1a ;
            rom[315] = 8'h21 ;
            rom[316] = 8'h2a ;
            rom[317] = 8'h3d ;
            rom[318] = 8'h17 ;
            rom[319] = 8'h02 ;
            rom[320] = 8'h32 ;
            rom[321] = 8'hea ;
            rom[322] = 8'h6b ;
            rom[323] = 8'h9a ;
            rom[324] = 8'hd6 ;
            rom[325] = 8'hab ;
            rom[326] = 8'h18 ;
            rom[327] = 8'hf1 ;
            rom[328] = 8'he5 ;
            rom[329] = 8'hdf ;
            rom[330] = 8'h05 ;
            rom[331] = 8'h2a ;
            rom[332] = 8'h28 ;
            rom[333] = 8'h25 ;
            rom[334] = 8'h10 ;
            rom[335] = 8'hc4 ;
            rom[336] = 8'h3b ;
            rom[337] = 8'hf4 ;
            rom[338] = 8'he6 ;
            rom[339] = 8'hff ;
            rom[340] = 8'hff ;
            rom[341] = 8'h2c ;
            rom[342] = 8'h2c ;
            rom[343] = 8'h41 ;
            rom[344] = 8'h03 ;
            rom[345] = 8'hc8 ;
            rom[346] = 8'h18 ;
            rom[347] = 8'h1b ;
            rom[348] = 8'hc9 ;
            rom[349] = 8'h1d ;
            rom[350] = 8'h21 ;
            rom[351] = 8'h30 ;
            rom[352] = 8'h2e ;
            rom[353] = 8'he2 ;
            rom[354] = 8'h5f ;
            rom[355] = 8'hc7 ;
            rom[356] = 8'hf3 ;
            rom[357] = 8'he7 ;
            rom[358] = 8'hee ;
            rom[359] = 8'h3a ;
            rom[360] = 8'hef ;
            rom[361] = 8'ha6 ;
            rom[362] = 8'h31 ;
            rom[363] = 8'hd0 ;
            rom[364] = 8'h31 ;
            rom[365] = 8'h23 ;
            rom[366] = 8'he5 ;
            rom[367] = 8'h10 ;
            rom[368] = 8'h1a ;
            rom[369] = 8'h5a ;
            rom[370] = 8'hdc ;
            rom[371] = 8'h07 ;
            rom[372] = 8'hf5 ;
            rom[373] = 8'h37 ;
            rom[374] = 8'h2c ;
            rom[375] = 8'he6 ;
            rom[376] = 8'h01 ;
            rom[377] = 8'h14 ;
            rom[378] = 8'h1b ;
            rom[379] = 8'hf0 ;
            rom[380] = 8'h1b ;
            rom[381] = 8'hf4 ;
            rom[382] = 8'he3 ;
            rom[383] = 8'hd0 ;
            rom[384] = 8'hd5 ;
            rom[385] = 8'hdf ;
            rom[386] = 8'h02 ;
            rom[387] = 8'h48 ;
            rom[388] = 8'hee ;
            rom[389] = 8'hee ;
            rom[390] = 8'hdb ;
            rom[391] = 8'hfa ;
            rom[392] = 8'he0 ;
            rom[393] = 8'h37 ;
            rom[394] = 8'h00 ;
            rom[395] = 8'hbd ;
            rom[396] = 8'h45 ;
            rom[397] = 8'hc6 ;
            rom[398] = 8'hed ;
            rom[399] = 8'h00 ;
            rom[400] = 8'hfa ;
            rom[401] = 8'hc2 ;
            rom[402] = 8'hf2 ;
            rom[403] = 8'h07 ;
            rom[404] = 8'hfe ;
            rom[405] = 8'hda ;
            rom[406] = 8'h00 ;
            rom[407] = 8'hd3 ;
            rom[408] = 8'h44 ;
            rom[409] = 8'h23 ;
            rom[410] = 8'hf4 ;
            rom[411] = 8'he7 ;
            rom[412] = 8'h53 ;
            rom[413] = 8'h01 ;
            rom[414] = 8'he5 ;
            rom[415] = 8'h17 ;
            rom[416] = 8'he6 ;
            rom[417] = 8'he1 ;
            rom[418] = 8'hcb ;
            rom[419] = 8'hff ;
            rom[420] = 8'hba ;
            rom[421] = 8'h19 ;
            rom[422] = 8'h1a ;
            rom[423] = 8'hfe ;
            rom[424] = 8'he1 ;
            rom[425] = 8'hec ;
            rom[426] = 8'he7 ;
            rom[427] = 8'h21 ;
            rom[428] = 8'h43 ;
            rom[429] = 8'h22 ;
            rom[430] = 8'hdf ;
            rom[431] = 8'hed ;
            rom[432] = 8'h17 ;
            rom[433] = 8'he2 ;
            rom[434] = 8'hcc ;
            rom[435] = 8'hf2 ;
            rom[436] = 8'h1a ;
            rom[437] = 8'hab ;
            rom[438] = 8'hfc ;
            rom[439] = 8'h01 ;
            rom[440] = 8'h10 ;
            rom[441] = 8'h00 ;
            rom[442] = 8'hcc ;
            rom[443] = 8'hac ;
            rom[444] = 8'h15 ;
            rom[445] = 8'h28 ;
            rom[446] = 8'h0b ;
            rom[447] = 8'h58 ;
            rom[448] = 8'hfd ;
            rom[449] = 8'hdf ;
            rom[450] = 8'he0 ;
            rom[451] = 8'hf1 ;
            rom[452] = 8'hbb ;
            rom[453] = 8'hfc ;
            rom[454] = 8'h1f ;
            rom[455] = 8'h11 ;
            rom[456] = 8'hdc ;
            rom[457] = 8'he1 ;
            rom[458] = 8'he1 ;
            rom[459] = 8'hbc ;
            rom[460] = 8'h1f ;
            rom[461] = 8'h52 ;
            rom[462] = 8'h03 ;
            rom[463] = 8'h0b ;
            rom[464] = 8'hdf ;
            rom[465] = 8'hfc ;
            rom[466] = 8'hfd ;
            rom[467] = 8'he7 ;
            rom[468] = 8'h02 ;
            rom[469] = 8'hcb ;
            rom[470] = 8'hd4 ;
            rom[471] = 8'ha9 ;
            rom[472] = 8'h37 ;
            rom[473] = 8'he8 ;
            rom[474] = 8'hdc ;
            rom[475] = 8'hc7 ;
            rom[476] = 8'h36 ;
            rom[477] = 8'h00 ;
            rom[478] = 8'hd0 ;
            rom[479] = 8'h3b ;
            rom[480] = 8'hec ;
            rom[481] = 8'he3 ;
            rom[482] = 8'h03 ;
            rom[483] = 8'h27 ;
            rom[484] = 8'h1d ;
            rom[485] = 8'hfe ;
            rom[486] = 8'h35 ;
            rom[487] = 8'h2e ;
            rom[488] = 8'hd7 ;
            rom[489] = 8'h12 ;
            rom[490] = 8'he9 ;
            rom[491] = 8'hc0 ;
            rom[492] = 8'h12 ;
            rom[493] = 8'hdd ;
            rom[494] = 8'hea ;
            rom[495] = 8'hd9 ;
            rom[496] = 8'hd5 ;
            rom[497] = 8'h03 ;
            rom[498] = 8'hde ;
            rom[499] = 8'hb7 ;
            rom[500] = 8'h36 ;
            rom[501] = 8'hf3 ;
            rom[502] = 8'h0d ;
            rom[503] = 8'he1 ;
            rom[504] = 8'h09 ;
            rom[505] = 8'hf6 ;
            rom[506] = 8'h1d ;
            rom[507] = 8'he9 ;
            rom[508] = 8'hdd ;
            rom[509] = 8'h13 ;
            rom[510] = 8'h2e ;
            rom[511] = 8'he7 ;
            rom[512] = 8'h18 ;
            rom[513] = 8'hd7 ;
            rom[514] = 8'hf0 ;
            rom[515] = 8'h42 ;
            rom[516] = 8'h0b ;
            rom[517] = 8'hc3 ;
            rom[518] = 8'h29 ;
            rom[519] = 8'h2a ;
            rom[520] = 8'hfb ;
            rom[521] = 8'he9 ;
            rom[522] = 8'he6 ;
            rom[523] = 8'h1d ;
            rom[524] = 8'hc8 ;
            rom[525] = 8'h11 ;
            rom[526] = 8'hee ;
            rom[527] = 8'hf2 ;
            rom[528] = 8'h0a ;
            rom[529] = 8'h2e ;
            rom[530] = 8'had ;
            rom[531] = 8'hbe ;
            rom[532] = 8'h0f ;
            rom[533] = 8'h02 ;
            rom[534] = 8'hd3 ;
            rom[535] = 8'hde ;
            rom[536] = 8'hdc ;
            rom[537] = 8'hd0 ;
            rom[538] = 8'hc9 ;
            rom[539] = 8'hf6 ;
            rom[540] = 8'he0 ;
            rom[541] = 8'h2a ;
            rom[542] = 8'h17 ;
            rom[543] = 8'hf3 ;
            rom[544] = 8'hff ;
            rom[545] = 8'h25 ;
            rom[546] = 8'h0e ;
            rom[547] = 8'h0b ;
            rom[548] = 8'hec ;
            rom[549] = 8'hfc ;
            rom[550] = 8'h47 ;
            rom[551] = 8'hf5 ;
            rom[552] = 8'h20 ;
            rom[553] = 8'hc6 ;
            rom[554] = 8'h05 ;
            rom[555] = 8'h01 ;
            rom[556] = 8'hc5 ;
            rom[557] = 8'h42 ;
            rom[558] = 8'hfb ;
            rom[559] = 8'hf7 ;
            rom[560] = 8'h35 ;
            rom[561] = 8'hdd ;
            rom[562] = 8'he9 ;
            rom[563] = 8'hab ;
            rom[564] = 8'h25 ;
            rom[565] = 8'hde ;
            rom[566] = 8'hc5 ;
            rom[567] = 8'hbb ;
            rom[568] = 8'hf0 ;
            rom[569] = 8'hce ;
            rom[570] = 8'hed ;
            rom[571] = 8'h0f ;
            rom[572] = 8'hf8 ;
            rom[573] = 8'hed ;
            rom[574] = 8'h1e ;
            rom[575] = 8'hd0 ;
            rom[576] = 8'he7 ;
            rom[577] = 8'h01 ;
            rom[578] = 8'h07 ;
            rom[579] = 8'hcd ;
            rom[580] = 8'h0f ;
            rom[581] = 8'hf8 ;
            rom[582] = 8'hb9 ;
            rom[583] = 8'hb9 ;
            rom[584] = 8'hd4 ;
            rom[585] = 8'h8c ;
            rom[586] = 8'h33 ;
            rom[587] = 8'h19 ;
            rom[588] = 8'hff ;
            rom[589] = 8'hf1 ;
            rom[590] = 8'hda ;
            rom[591] = 8'h19 ;
            rom[592] = 8'h1e ;
            rom[593] = 8'hf9 ;
            rom[594] = 8'hec ;
            rom[595] = 8'h09 ;
            rom[596] = 8'hf8 ;
            rom[597] = 8'hfc ;
            rom[598] = 8'h18 ;
            rom[599] = 8'hf7 ;
            rom[600] = 8'hee ;
            rom[601] = 8'hfe ;
            rom[602] = 8'hb4 ;
            rom[603] = 8'hf3 ;
            rom[604] = 8'h0b ;
            rom[605] = 8'h2e ;
            rom[606] = 8'hf5 ;
            rom[607] = 8'hfe ;
            rom[608] = 8'hbe ;
            rom[609] = 8'h14 ;
            rom[610] = 8'h1e ;
            rom[611] = 8'hd9 ;
            rom[612] = 8'hfd ;
            rom[613] = 8'h1a ;
            rom[614] = 8'h17 ;
            rom[615] = 8'h0e ;
            rom[616] = 8'hf2 ;
            rom[617] = 8'hc5 ;
            rom[618] = 8'h2a ;
            rom[619] = 8'h09 ;
            rom[620] = 8'h2c ;
            rom[621] = 8'h18 ;
            rom[622] = 8'h03 ;
            rom[623] = 8'hbc ;
            rom[624] = 8'h25 ;
            rom[625] = 8'h02 ;
            rom[626] = 8'hef ;
            rom[627] = 8'h1b ;
            rom[628] = 8'hd9 ;
            rom[629] = 8'hfb ;
            rom[630] = 8'h22 ;
            rom[631] = 8'hff ;
            rom[632] = 8'hd7 ;
            rom[633] = 8'hc7 ;
            rom[634] = 8'h17 ;
            rom[635] = 8'hf3 ;
            rom[636] = 8'he0 ;
            rom[637] = 8'h16 ;
            rom[638] = 8'h06 ;
            rom[639] = 8'h0c ;
            rom[640] = 8'hd7 ;
            rom[641] = 8'he7 ;
            rom[642] = 8'h33 ;
            rom[643] = 8'h2e ;
            rom[644] = 8'hc8 ;
            rom[645] = 8'h0e ;
            rom[646] = 8'he5 ;
            rom[647] = 8'h2e ;
            rom[648] = 8'h0a ;
            rom[649] = 8'ha9 ;
            rom[650] = 8'h2b ;
            rom[651] = 8'hf6 ;
            rom[652] = 8'h23 ;
            rom[653] = 8'he2 ;
            rom[654] = 8'h24 ;
            rom[655] = 8'hba ;
            rom[656] = 8'hda ;
            rom[657] = 8'h25 ;
            rom[658] = 8'hea ;
            rom[659] = 8'hfe ;
            rom[660] = 8'h28 ;
            rom[661] = 8'h36 ;
            rom[662] = 8'h3f ;
            rom[663] = 8'h02 ;
            rom[664] = 8'hae ;
            rom[665] = 8'heb ;
            rom[666] = 8'h08 ;
            rom[667] = 8'h1a ;
            rom[668] = 8'h08 ;
            rom[669] = 8'ha5 ;
            rom[670] = 8'h13 ;
            rom[671] = 8'h07 ;
            rom[672] = 8'hcb ;
            rom[673] = 8'h03 ;
            rom[674] = 8'h05 ;
            rom[675] = 8'h00 ;
            rom[676] = 8'hf1 ;
            rom[677] = 8'hd1 ;
            rom[678] = 8'hba ;
            rom[679] = 8'hda ;
            rom[680] = 8'he8 ;
            rom[681] = 8'h2d ;
            rom[682] = 8'hd5 ;
            rom[683] = 8'h2c ;
            rom[684] = 8'he9 ;
            rom[685] = 8'hb4 ;
            rom[686] = 8'h07 ;
            rom[687] = 8'hee ;
            rom[688] = 8'hc2 ;
            rom[689] = 8'h05 ;
            rom[690] = 8'hf5 ;
            rom[691] = 8'h21 ;
            rom[692] = 8'h14 ;
            rom[693] = 8'hfe ;
            rom[694] = 8'h27 ;
            rom[695] = 8'h1b ;
            rom[696] = 8'h55 ;
            rom[697] = 8'he5 ;
            rom[698] = 8'hda ;
            rom[699] = 8'hd3 ;
            rom[700] = 8'hda ;
            rom[701] = 8'h35 ;
            rom[702] = 8'hdb ;
            rom[703] = 8'hc8 ;
            rom[704] = 8'he3 ;
            rom[705] = 8'hdf ;
            rom[706] = 8'he8 ;
            rom[707] = 8'h32 ;
            rom[708] = 8'hac ;
            rom[709] = 8'he3 ;
            rom[710] = 8'he1 ;
            rom[711] = 8'h28 ;
            rom[712] = 8'hf6 ;
            rom[713] = 8'hea ;
            rom[714] = 8'hc8 ;
            rom[715] = 8'h51 ;
            rom[716] = 8'he4 ;
            rom[717] = 8'h05 ;
            rom[718] = 8'hf8 ;
            rom[719] = 8'h17 ;
            rom[720] = 8'hc3 ;
            rom[721] = 8'hfa ;
            rom[722] = 8'hc4 ;
            rom[723] = 8'h1b ;
            rom[724] = 8'he2 ;
            rom[725] = 8'hb7 ;
            rom[726] = 8'he6 ;
            rom[727] = 8'h0c ;
            rom[728] = 8'h0b ;
            rom[729] = 8'hc7 ;
            rom[730] = 8'hde ;
            rom[731] = 8'h00 ;
            rom[732] = 8'h25 ;
            rom[733] = 8'h25 ;
            rom[734] = 8'hc9 ;
            rom[735] = 8'h21 ;
            rom[736] = 8'h18 ;
            rom[737] = 8'h05 ;
            rom[738] = 8'h0a ;
            rom[739] = 8'h09 ;
            rom[740] = 8'hdc ;
            rom[741] = 8'hbd ;
            rom[742] = 8'hcf ;
            rom[743] = 8'hf3 ;
            rom[744] = 8'hf5 ;
            rom[745] = 8'hf6 ;
            rom[746] = 8'hee ;
            rom[747] = 8'h43 ;
            rom[748] = 8'hbc ;
            rom[749] = 8'he7 ;
            rom[750] = 8'hfe ;
            rom[751] = 8'hf1 ;
            rom[752] = 8'h12 ;
            rom[753] = 8'he3 ;
            rom[754] = 8'h23 ;
            rom[755] = 8'h4f ;
            rom[756] = 8'hef ;
            rom[757] = 8'hea ;
            rom[758] = 8'hee ;
            rom[759] = 8'hde ;
            rom[760] = 8'h17 ;
            rom[761] = 8'he1 ;
            rom[762] = 8'h17 ;
            rom[763] = 8'h03 ;
            rom[764] = 8'h3e ;
            rom[765] = 8'hed ;
            rom[766] = 8'hfe ;
            rom[767] = 8'he3 ;
            rom[768] = 8'hef ;
            rom[769] = 8'h0b ;
            rom[770] = 8'hf3 ;
            rom[771] = 8'hc3 ;
            rom[772] = 8'hf9 ;
            rom[773] = 8'h20 ;
            rom[774] = 8'h06 ;
            rom[775] = 8'hff ;
            rom[776] = 8'he1 ;
            rom[777] = 8'h08 ;
            rom[778] = 8'hf5 ;
            rom[779] = 8'he7 ;
            rom[780] = 8'h22 ;
            rom[781] = 8'he3 ;
            rom[782] = 8'hdf ;
            rom[783] = 8'hd9 ;
            rom[784] = 8'hf1 ;
            rom[785] = 8'he8 ;
            rom[786] = 8'hc8 ;
            rom[787] = 8'hcd ;
            rom[788] = 8'hf3 ;
            rom[789] = 8'h17 ;
            rom[790] = 8'hd5 ;
            rom[791] = 8'h37 ;
            rom[792] = 8'h40 ;
            rom[793] = 8'hd9 ;
            rom[794] = 8'h51 ;
            rom[795] = 8'hc2 ;
            rom[796] = 8'hd4 ;
            rom[797] = 8'h12 ;
            rom[798] = 8'h34 ;
            rom[799] = 8'hed ;
            rom[800] = 8'h38 ;
            rom[801] = 8'h14 ;
            rom[802] = 8'hcb ;
            rom[803] = 8'hfb ;
            rom[804] = 8'hc7 ;
            rom[805] = 8'h2c ;
            rom[806] = 8'hdb ;
            rom[807] = 8'h1f ;
            rom[808] = 8'h18 ;
            rom[809] = 8'h10 ;
            rom[810] = 8'hd8 ;
            rom[811] = 8'h32 ;
            rom[812] = 8'he2 ;
            rom[813] = 8'h00 ;
            rom[814] = 8'hdd ;
            rom[815] = 8'h3c ;
            rom[816] = 8'he2 ;
            rom[817] = 8'h30 ;
            rom[818] = 8'hef ;
            rom[819] = 8'hf8 ;
            rom[820] = 8'h2c ;
            rom[821] = 8'h16 ;
            rom[822] = 8'hba ;
            rom[823] = 8'h40 ;
            rom[824] = 8'he2 ;
            rom[825] = 8'hed ;
            rom[826] = 8'h08 ;
            rom[827] = 8'hbc ;
            rom[828] = 8'h0a ;
            rom[829] = 8'hff ;
            rom[830] = 8'h37 ;
            rom[831] = 8'hd7 ;
            rom[832] = 8'h4b ;
            rom[833] = 8'heb ;
            rom[834] = 8'hb3 ;
            rom[835] = 8'h2c ;
            rom[836] = 8'h0c ;
            rom[837] = 8'h0c ;
            rom[838] = 8'he7 ;
            rom[839] = 8'h05 ;
            rom[840] = 8'hee ;
            rom[841] = 8'he1 ;
            rom[842] = 8'he1 ;
            rom[843] = 8'he3 ;
            rom[844] = 8'hc0 ;
            rom[845] = 8'h1b ;
            rom[846] = 8'h15 ;
            rom[847] = 8'h29 ;
            rom[848] = 8'h55 ;
            rom[849] = 8'he8 ;
            rom[850] = 8'he9 ;
            rom[851] = 8'h38 ;
            rom[852] = 8'h05 ;
            rom[853] = 8'hdd ;
            rom[854] = 8'hd2 ;
            rom[855] = 8'h3a ;
            rom[856] = 8'hde ;
            rom[857] = 8'h0b ;
            rom[858] = 8'h3b ;
            rom[859] = 8'hd0 ;
            rom[860] = 8'hfa ;
            rom[861] = 8'hba ;
            rom[862] = 8'h28 ;
            rom[863] = 8'hb4 ;
        end
    always
        @(*)
        begin
            data = rom[addr] ;
        end
endmodule



